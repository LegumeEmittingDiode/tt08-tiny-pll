module tt08_integration (
	VGND,
	VPWR,
	clk_ref_0,
	clk_ref_1,
	clk_ref_2,
	clk_ref_3,
	div_fb0_0,
	div_fb0_1,
	div_fb0_2,
	div_fb0_3,
	div_fb1_0,
	div_fb1_1,
	div_fb1_2,
	div_fb1_3,
	div_fb2_0,
	div_fb2_1,
	div_fb2_2,
	div_fb2_3,
	div_fb3_0,
	div_fb3_1,
	div_fb3_2,
	div_fb3_3,
	div_out0_0,
	div_out0_1,
	div_out0_2,
	div_out0_3,
	div_out1_0,
	div_out1_1,
	div_out1_2,
	div_out1_3,
	div_out2_0,
	div_out2_1,
	div_out2_2,
	div_out2_3,
	div_out3_0,
	div_out3_1,
	div_out3_2,
	div_out3_3,
	enb_0,
	enb_1,
	enb_2,
	enb_3,
	clk_out_0,
	clk_out_1,
	clk_out_2,
	clk_out_3,
	adc_out
);

input VGND;
input VPWR;
input clk_ref_0;
input clk_ref_1;
input clk_ref_2;
input clk_ref_3;
input div_fb0_0;
input div_fb0_1;
input div_fb0_2;
input div_fb0_3;
input div_fb1_0;
input div_fb1_1;
input div_fb1_2;
input div_fb1_3;
input div_fb2_0;
input div_fb2_1;
input div_fb2_2;
input div_fb2_3;
input div_fb3_0;
input div_fb3_1;
input div_fb3_2;
input div_fb3_3;
input div_out0_0;
input div_out0_1;
input div_out0_2;
input div_out0_3;
input div_out1_0;
input div_out1_1;
input div_out1_2;
input div_out1_3;
input div_out2_0;
input div_out2_1;
input div_out2_2;
input div_out2_3;
input div_out3_0;
input div_out3_1;
input div_out3_2;
input div_out3_3;
input enb_0;
input enb_1;
input enb_2;
input enb_3;
output clk_out_0;
output clk_out_1;
output clk_out_2;
output clk_out_3;
output adc_out;

endmodule

