* NGSPICE file created from tt_um_tiny_pll.ext - technology: sky130A

.subckt sky130_fd_sc_hd__decap_6 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.97
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.97
.ends

.subckt sky130_fd_sc_hd__clkbuf_1 VGND VPWR VNB VPB X A
X0 VPWR a_75_212# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X1 a_75_212# A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2 a_75_212# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X3 VGND a_75_212# X VNB sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_3 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=0.59
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=0.59
.ends

.subckt sky130_fd_sc_hd__clkbuf_2 VGND VPWR VNB VPB A X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1625 pd=1.325 as=0.265 ps=2.53 w=1 l=0.15
X1 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.06825 pd=0.745 as=0.1113 ps=1.37 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.1625 ps=1.325 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.06825 ps=0.745 w=0.42 l=0.15
X5 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfrtp_1 VGND VPWR VNB VPB CLK D RESET_B Q
X0 a_805_47# a_761_289# a_639_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1 a_1217_47# a_27_47# a_1108_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2 a_1283_21# a_1108_47# a_1462_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X3 a_651_413# a_27_47# a_543_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X4 a_1108_47# a_193_47# a_761_289# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X5 VGND RESET_B a_805_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X6 Q a_1283_21# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X7 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_448_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 a_761_289# a_543_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X10 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 a_1108_47# a_27_47# a_761_289# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X12 a_1462_47# RESET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X13 a_543_47# a_27_47# a_448_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X14 a_543_47# a_193_47# a_448_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X15 a_448_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X16 VPWR a_1283_21# a_1270_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VPWR a_1108_47# a_1283_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 a_1270_413# a_193_47# a_1108_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X19 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 a_1283_21# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X21 VPWR a_761_289# a_651_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X22 Q a_1283_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X23 a_639_47# a_193_47# a_543_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X24 VGND a_1283_21# a_1217_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X25 a_651_413# RESET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X26 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 a_761_289# a_543_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
.ends

.subckt sky130_ef_sc_hd__decap_12 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=4.73
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=4.73
.ends

.subckt sky130_fd_sc_hd__mux2_1 VGND VPWR VNB VPB X A1 S A0
X0 VPWR a_505_21# a_535_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X1 a_505_21# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1176 pd=1.4 as=0.0693 ps=0.75 w=0.42 l=0.15
X2 a_218_374# S VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.15835 ps=1.395 w=0.42 l=0.15
X3 VGND a_505_21# a_439_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1449 pd=1.11 as=0.0693 ps=0.75 w=0.42 l=0.15
X4 a_76_199# A0 a_218_374# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1932 pd=1.34 as=0.07665 ps=0.785 w=0.42 l=0.15
X5 a_505_21# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1449 ps=1.11 w=0.42 l=0.15
X6 a_439_47# A0 a_76_199# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.09975 ps=0.895 w=0.42 l=0.15
X7 a_535_374# A1 a_76_199# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.1932 ps=1.34 w=0.42 l=0.15
X8 a_76_199# A1 a_218_47# VNB sky130_fd_pr__nfet_01v8 ad=0.09975 pd=0.895 as=0.0693 ps=0.75 w=0.42 l=0.15
X9 a_218_47# S VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.11285 ps=1.045 w=0.42 l=0.15
X10 VPWR a_76_199# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.15835 pd=1.395 as=0.26 ps=2.52 w=1 l=0.15
X11 VGND a_76_199# X VNB sky130_fd_pr__nfet_01v8 ad=0.11285 pd=1.045 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nand4b_1 VGND VPWR VNB VPB Y C B D A_N
X0 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.195 pd=1.39 as=0.1925 ps=1.385 w=1 l=0.15
X1 a_232_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.118125 ps=1.04 w=0.65 l=0.15
X2 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1925 pd=1.385 as=0.135 ps=1.27 w=1 l=0.15
X3 VPWR A_N a_41_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14575 pd=1.335 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VPWR a_41_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.195 ps=1.39 w=1 l=0.15
X5 a_316_47# C a_232_47# VNB sky130_fd_pr__nfet_01v8 ad=0.125125 pd=1.035 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 Y a_41_93# a_423_47# VNB sky130_fd_pr__nfet_01v8 ad=0.2275 pd=2 as=0.12675 ps=1.04 w=0.65 l=0.15
X7 a_423_47# B a_316_47# VNB sky130_fd_pr__nfet_01v8 ad=0.12675 pd=1.04 as=0.125125 ps=1.035 w=0.65 l=0.15
X8 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.14575 ps=1.335 w=1 l=0.15
X9 VGND A_N a_41_93# VNB sky130_fd_pr__nfet_01v8 ad=0.118125 pd=1.04 as=0.1113 ps=1.37 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dfstp_1 VPWR VGND VNB VPB Q SET_B D CLK
X0 VGND a_652_21# a_586_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0882 pd=0.84 as=0.06705 ps=0.75 w=0.42 l=0.15
X1 a_956_413# a_476_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0483 pd=0.65 as=0.0567 ps=0.69 w=0.42 l=0.15
X2 VPWR a_476_47# a_652_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X3 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X4 a_586_47# a_193_47# a_476_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.072 ps=0.76 w=0.36 l=0.15
X5 a_1056_47# a_476_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X6 a_476_47# a_27_47# a_381_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.0935 ps=0.965 w=0.36 l=0.15
X7 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12495 pd=1.175 as=0.2184 ps=2.2 w=0.84 l=0.15
X8 a_652_21# SET_B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0798 ps=0.8 w=0.42 l=0.15
X9 a_1224_47# a_27_47# a_1032_413# VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0693 ps=0.75 w=0.42 l=0.15
X10 a_562_413# a_27_47# a_476_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0945 pd=0.87 as=0.0567 ps=0.69 w=0.42 l=0.15
X11 VGND a_1032_413# a_1602_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X12 VPWR a_1182_261# a_1140_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X13 Q a_1602_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.149 ps=1.325 w=1 l=0.15
X14 a_1032_413# a_193_47# a_1056_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0693 pd=0.75 as=0.0441 ps=0.63 w=0.42 l=0.15
X15 a_476_47# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.12495 ps=1.175 w=0.42 l=0.15
X16 a_1296_47# a_1182_261# a_1224_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0483 pd=0.65 as=0.0441 ps=0.63 w=0.42 l=0.15
X17 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X18 VPWR a_652_21# a_562_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0798 pd=0.8 as=0.0945 ps=0.87 w=0.42 l=0.15
X19 VPWR SET_B a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.12285 pd=1.17 as=0.1092 ps=1.36 w=0.42 l=0.15
X20 a_1032_413# a_27_47# a_956_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0483 ps=0.65 w=0.42 l=0.15
X21 a_1182_261# a_1032_413# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12285 ps=1.17 w=0.84 l=0.15
X22 Q a_1602_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X23 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X24 a_1140_413# a_193_47# a_1032_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0441 pd=0.63 as=0.0819 ps=0.81 w=0.42 l=0.15
X25 VPWR a_1032_413# a_1602_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X26 a_796_47# SET_B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.0882 ps=0.84 w=0.42 l=0.15
X27 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0935 pd=0.965 as=0.1664 ps=1.8 w=0.64 l=0.15
X28 a_1182_261# a_1032_413# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1404 pd=1.6 as=0.1137 ps=1.01 w=0.54 l=0.15
X29 a_652_21# a_476_47# a_796_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X30 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X31 VGND SET_B a_1296_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1137 pd=1.01 as=0.0483 ps=0.65 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__decap_4 VGND VPWR VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=1.05
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=1.05
.ends

.subckt sky130_fd_sc_hd__clkbuf_4 VGND VPWR VNB VPB A X
X0 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.265 ps=2.53 w=1 l=0.15
X1 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.1218 pd=1.42 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.0588 ps=0.7 w=0.42 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.07035 pd=0.755 as=0.1113 ps=1.37 w=0.42 l=0.15
X6 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.14 ps=1.28 w=1 l=0.15
X7 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.07035 ps=0.755 w=0.42 l=0.15
X8 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.165 ps=1.33 w=1 l=0.15
X9 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14 pd=1.28 as=0.14 ps=1.28 w=1 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4bb_2 VGND VPWR VNB VPB Y B A D_N C_N
X0 Y a_27_410# a_336_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 a_336_297# a_201_93# a_418_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 Y a_201_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.221 ps=1.98 w=0.65 l=0.15
X4 Y a_27_410# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X6 a_418_297# a_201_93# a_336_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X7 VGND D_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 VPWR D_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X9 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.17875 pd=1.85 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_776_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.275 pd=2.55 as=0.135 ps=1.27 w=1 l=0.15
X12 a_201_93# C_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1226 ps=1.32 w=0.42 l=0.15
X13 a_201_93# C_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X14 VPWR A a_776_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X15 a_776_297# B a_418_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X16 VGND a_201_93# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 a_336_297# a_27_410# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X18 a_418_297# B a_776_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X19 VGND a_27_410# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_4 VPWR VGND VNB VPB A X
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X3 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X9 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__buf_2 VPWR VGND VNB VPB X A
X0 VPWR a_27_47# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.265 pd=2.53 as=0.135 ps=1.27 w=1 l=0.15
X1 X a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.149 ps=1.325 w=1 l=0.15
X2 VPWR A a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.149 pd=1.325 as=0.1664 ps=1.8 w=0.64 l=0.15
X3 X a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.097 ps=0.975 w=0.65 l=0.15
X4 VGND a_27_47# X VNB sky130_fd_pr__nfet_01v8 ad=0.17225 pd=1.83 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 VGND A a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__dlymetal6s2s_1 VPWR VGND VNB VPB X A
X0 a_558_47# a_381_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1 VGND X a_381_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 a_841_47# a_664_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X3 VPWR A a_62_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X4 VGND A a_62_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_558_47# a_381_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X6 X a_62_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X7 VPWR X a_381_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X8 a_841_47# a_664_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X9 X a_62_47# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X10 VPWR a_558_47# a_664_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 VGND a_558_47# a_664_47# VNB sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__and4bb_1 VGND VPWR VNB VPB A_N B_N C D X
X0 VPWR D a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.172 pd=1.46 as=0.0777 ps=0.79 w=0.42 l=0.15
X1 a_223_47# B_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1386 pd=1.5 as=0.0588 ps=0.7 w=0.42 l=0.15
X2 a_515_93# a_223_47# a_429_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
X3 a_223_47# B_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1344 pd=1.48 as=0.0588 ps=0.7 w=0.42 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X5 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.168 ps=1.64 w=0.42 l=0.15
X6 X a_343_93# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.172 ps=1.46 w=1 l=0.15
X7 a_429_93# a_27_47# a_343_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0588 pd=0.7 as=0.1176 ps=1.4 w=0.42 l=0.15
X8 VGND D a_615_93# VNB sky130_fd_pr__nfet_01v8 ad=0.1265 pd=1.11 as=0.0777 ps=0.79 w=0.42 l=0.15
X9 a_343_93# C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X10 a_343_93# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.1218 ps=1.42 w=0.42 l=0.15
X11 a_615_93# C a_515_93# VNB sky130_fd_pr__nfet_01v8 ad=0.0777 pd=0.79 as=0.0735 ps=0.77 w=0.42 l=0.15
X12 X a_343_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1654 pd=1.82 as=0.1265 ps=1.11 w=0.65 l=0.15
X13 VPWR a_223_47# a_343_93# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0735 pd=0.77 as=0.0588 ps=0.7 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__conb_1 VGND VPWR VNB VPB LO HI
X0 VPWR HI sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1 LO VGND sky130_fd_pr__res_generic_po w=0.48 l=0.045
.ends

.subckt sky130_fd_sc_hd__decap_8 VPWR VGND VNB VPB
X0 VPWR VGND VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0.4524 ps=4.52 w=0.87 l=2.89
X1 VGND VPWR VGND VNB sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0.286 ps=3.24 w=0.55 l=2.89
.ends

.subckt sky130_fd_sc_hd__nand4b_2 VGND VPWR VNB VPB A_N Y B C D
X0 Y a_27_47# a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1 a_465_47# B a_215_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND D a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.117 ps=1.01 w=0.65 l=0.15
X3 a_215_47# B a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR A_N a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_655_47# D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 a_655_47# C a_465_47# VNB sky130_fd_pr__nfet_01v8 ad=0.117 pd=1.01 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 VPWR B Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.37 pd=1.74 as=0.135 ps=1.27 w=1 l=0.15
X8 Y B VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X9 a_465_47# C a_655_47# VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X10 VPWR a_27_47# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 VPWR C Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.18 pd=1.36 as=0.135 ps=1.27 w=1 l=0.15
X12 VPWR D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.4 pd=2.8 as=0.135 ps=1.27 w=1 l=0.15
X13 Y D VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.18 ps=1.36 w=1 l=0.15
X14 a_215_47# a_27_47# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 Y a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X16 Y C VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.37 ps=1.74 w=1 l=0.15
X17 VGND A_N a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4b_4 VGND VPWR VNB VPB B D_N A C Y
X0 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND D_N a_1191_21# VNB sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.169 ps=1.82 w=0.65 l=0.15
X3 a_803_297# a_1191_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X4 a_445_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y a_1191_21# a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X7 a_803_297# a_1191_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X10 Y a_1191_21# a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X11 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X12 Y a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X14 VPWR D_N a_1191_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.28 pd=2.56 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X17 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X18 a_27_297# B a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X19 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 VGND a_1191_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X21 VGND a_1191_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X22 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 a_445_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X25 a_803_297# C a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X26 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X27 a_27_297# B a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X28 a_445_297# C a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 a_803_297# C a_445_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 Y a_1191_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X31 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X32 a_445_297# C a_803_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4b_2 VGND VPWR VNB VPB A B C Y D_N
X0 VPWR D_N a_694_21# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X1 a_27_297# B a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2 a_474_297# a_694_21# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X3 a_277_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 Y a_694_21# a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X6 VGND D_N a_694_21# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.1092 ps=1.36 w=0.42 l=0.15
X7 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X8 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X9 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X11 a_474_297# C a_277_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X12 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X13 Y a_694_21# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_277_297# C a_474_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X15 VGND a_694_21# Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X17 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4bb_1 VGND VPWR VNB VPB A Y B D_N C_N
X0 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10725 ps=0.98 w=0.65 l=0.15
X1 VGND a_27_410# Y VNB sky130_fd_pr__nfet_01v8 ad=0.10725 pd=0.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X2 VGND C_N a_27_410# VNB sky130_fd_pr__nfet_01v8 ad=0.0609 pd=0.71 as=0.1092 ps=1.36 w=0.42 l=0.15
X3 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 VPWR C_N a_27_410# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1226 pd=1.32 as=0.1092 ps=1.36 w=0.42 l=0.15
X5 a_205_93# D_N VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0609 ps=0.71 w=0.42 l=0.15
X6 VPWR A a_573_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X7 a_205_93# D_N VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1085 pd=1.36 as=0.1226 ps=1.32 w=0.42 l=0.15
X8 a_477_297# a_27_410# a_393_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.165 pd=1.33 as=0.135 ps=1.27 w=1 l=0.15
X9 a_573_297# B a_477_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.165 ps=1.33 w=1 l=0.15
X10 a_393_297# a_205_93# Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.2559 ps=2.52 w=1 l=0.15
X11 Y a_205_93# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
.ends

.subckt sky130_fd_sc_hd__mux4_2 VGND VPWR VNB VPB S0 A2 A3 S1 A1 A0 X
X0 a_600_345# S1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_788_316# S1 a_288_47# VNB sky130_fd_pr__nfet_01v8 ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2 VPWR A3 a_372_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1645 ps=1.33 w=0.64 l=0.15
X3 a_872_316# a_600_345# a_788_316# VNB sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X4 VPWR S0 a_27_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X5 a_1279_413# S0 a_872_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.10535 pd=0.995 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 VGND a_788_316# X VNB sky130_fd_pr__nfet_01v8 ad=0.221 pd=1.98 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_1060_369# A1 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.13775 pd=1.165 as=0.1664 ps=1.8 w=0.64 l=0.15
X8 a_872_316# a_27_47# a_1060_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.13775 ps=1.165 w=0.42 l=0.15
X9 a_193_47# A2 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.0567 ps=0.69 w=0.42 l=0.15
X10 a_1064_47# A1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.0786 pd=0.805 as=0.1092 ps=1.36 w=0.42 l=0.15
X11 a_1281_47# a_27_47# a_872_316# VNB sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.072 ps=0.76 w=0.36 l=0.15
X12 a_872_316# S1 a_788_316# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1404 pd=1.6 as=0.0729 ps=0.81 w=0.54 l=0.15
X13 a_872_316# S0 a_1064_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.072 pd=0.76 as=0.0786 ps=0.805 w=0.36 l=0.15
X14 X a_788_316# VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.10675 ps=1.005 w=0.65 l=0.15
X15 a_788_316# a_600_345# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0729 pd=0.81 as=0.1404 ps=1.6 w=0.54 l=0.15
X16 a_372_413# a_27_47# a_288_47# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1645 pd=1.33 as=0.0567 ps=0.69 w=0.42 l=0.15
X17 VGND A3 a_397_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0819 pd=0.81 as=0.06705 ps=0.75 w=0.42 l=0.15
X18 a_600_345# S1 VGND VNB sky130_fd_pr__nfet_01v8 ad=0.1134 pd=1.38 as=0.0819 ps=0.81 w=0.42 l=0.15
X19 a_193_369# A2 VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.09575 pd=0.965 as=0.0864 ps=0.91 w=0.64 l=0.15
X20 VPWR a_788_316# X VPB sky130_fd_pr__pfet_01v8_hvt ad=0.34 pd=2.68 as=0.135 ps=1.27 w=1 l=0.15
X21 a_288_47# S0 a_193_369# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.09575 ps=0.965 w=0.42 l=0.15
X22 VGND A0 a_1281_47# VNB sky130_fd_pr__nfet_01v8 ad=0.10675 pd=1.005 as=0.066 ps=0.745 w=0.42 l=0.15
X23 a_397_47# S0 a_288_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.06705 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X24 X a_788_316# VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.154 ps=1.335 w=1 l=0.15
X25 a_288_47# a_27_47# a_193_47# VNB sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.066 ps=0.745 w=0.36 l=0.15
X26 VGND S0 a_27_47# VNB sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VPWR A0 a_1279_413# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.10535 ps=0.995 w=0.64 l=0.15
.ends

.subckt sky130_fd_sc_hd__nor4_4 VGND VPWR VNB VPB A B Y D C
X0 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X4 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X5 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X6 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X8 Y C VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25675 ps=1.44 w=0.65 l=0.15
X9 Y D VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X10 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X11 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X12 Y A VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.182 ps=1.86 w=0.65 l=0.15
X13 VGND A Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X15 VGND B Y VNB sky130_fd_pr__nfet_01v8 ad=0.25675 pd=1.44 as=0.08775 ps=0.92 w=0.65 l=0.15
X16 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X17 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X18 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X19 VGND D Y VNB sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X20 a_807_297# C a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X21 VPWR A a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.28 ps=2.56 w=1 l=0.15
X22 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X23 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X24 Y B VGND VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X25 a_449_297# C a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X26 a_27_297# B a_449_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X27 a_807_297# D Y VPB sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X28 a_449_297# B a_27_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X29 Y D a_807_297# VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X30 a_27_297# A VPWR VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X31 VGND C Y VNB sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
.ends

.subckt tt08_integration div_fb0_1 div_fb1_1 div_fb2_1 div_fb3_1 div_out0_1 div_out2_1
+ div_out1_1 div_out3_1 div_out3_2 div_out1_2 div_out2_2 div_out0_2 div_fb3_2 div_fb2_2
+ div_fb1_2 div_fb0_2 div_out3_3 div_out1_3 div_out2_3 div_out0_3 div_fb3_3 div_fb2_3
+ div_fb1_3 div_fb0_3 div_fb0_0 div_fb1_0 div_fb2_0 div_fb3_0 div_out0_0 div_out2_0
+ div_out1_0 div_out3_0 enb_0 clk_ref_0 w_62_6889# w_62_2537# a_3660_7915# a_209_147#
+ w_62_10153# a_12261_8673# w_62_5801# a_3519_9941# a_13743_5587# a_127_7559# a_15289_9939#
+ a_127_3207# w_62_14505# a_15289_10483# w_62_7977# a_127_4295# w_62_3625# a_15289_2323#
+ w_62_9065# w_62_361# w_62_15593# w_62_11241# a_13661_5587# w_62_12329# a_3519_10499#
+ w_62_1449# a_11774_6622# a_3519_15381# a_127_5383# w_62_4713# a_3660_13355# a_15289_15379#
+ a_3660_12891# w_62_13417# a_12261_11891# a_12261_14113# a_6055_3079# a_209_11027#
+ a_14203_3207#
X0 w_62_14505# a_179_14265# a_127_14291# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X1 w_62_12329# a_11296_11803# a_11903_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2 a_12695_2157# a_12179_1785# a_12600_2145# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X3 w_62_10153# div_out0_2 a_13281_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X4 a_127_3207# a_13835_147# a_14079_665# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X5 a_12528_8129# a_12498_8015# a_12231_7737# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X6 a_1397_1235# div_fb0_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X7 a_3250_12481# a_2754_12267# a_3079_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X8 a_127_3207# clk_ref_0 a_3465_2351# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X9 a_127_3207# a_7331_4818# a_8109_7110# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X10 a_5225_1645# a_4971_332# a_4971_332# w_62_1449# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1 as=0.15 ps=1.6 w=0.5 l=0.15
X11 a_15126_8129# a_14407_7905# a_14563_8000# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X12 w_62_3625# a_127_3207# w_62_3625# w_62_3625# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=3.6192 ps=36.16 w=0.87 l=1.05
X13 a_127_3207# a_13835_13203# a_14079_13721# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X14 a_3379_15407# a_1225_15531# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X15 a_534_9031# a_1383_9699# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X16 a_127_3207# a_179_13177# a_127_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X17 a_13422_8307# a_12179_8313# a_13260_8685# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X18 a_1147_9101# a_534_9031# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X19 a_643_12115# a_127_12115# a_548_12115# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X20 a_5929_2573# a_5419_2297# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X21 a_11296_1387# a_11658_1235# a_11300_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X22 a_127_3207# w_62_4713# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=202.2677 ps=1.81328k w=0.55 l=4.73
X23 a_14801_11937# a_12854_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X24 a_13435_11001# a_13260_11027# a_13614_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X25 a_1370_11393# a_127_11027# a_1208_11027# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X26 a_12345_12115# a_12179_12115# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X27 w_62_10153# a_12174_8539# a_12179_9401# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X28 w_62_10153# a_14239_10483# a_14407_10457# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X29 a_8199_4858# a_6485_5594# a_9567_4858# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=0.5
X30 a_14109_13747# a_13835_13203# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X31 w_62_12329# a_15188_12633# a_15126_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X32 a_12174_923# a_1225_2475# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X33 a_1317_2157# a_293_1785# a_1208_2157# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X34 a_127_3207# a_15188_8012# a_15126_8129# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X35 w_62_11241# a_5225_11511# a_5225_11511# w_62_11241# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.125 ps=1 w=0.5 l=0.15
X36 a_13449_14541# div_out0_3 w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X37 a_14806_11179# a_14755_12115# a_14932_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X38 a_350_7915# a_446_8015# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X39 a_4150_8648# a_4910_8536# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X40 a_4150_14088# a_4910_13976# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X41 a_12803_1779# a_12345_1785# a_12695_2157# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X42 a_9193_6328# a_6485_6328# a_8019_7110# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=0.5
X43 a_397_11937# a_350_11803# a_179_11545# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X44 a_12695_1069# a_12179_697# a_12600_1057# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X45 a_127_3207# w_62_5801# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X46 a_13614_8673# a_12854_9939# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X47 a_1208_1069# a_127_697# a_861_665# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X48 w_62_10153# a_1371_10457# a_122_11179# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X49 a_534_14471# a_1383_15139# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X50 a_13260_2157# a_12179_1785# a_12913_1753# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X51 a_13449_13203# div_out1_3 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X52 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X53 a_3140_9395# a_1783_8851# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X54 a_127_3207# a_4315_2297# a_3617_1387# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X55 a_485_2573# a_397_2475# a_403_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X56 a_13940_10861# a_13541_10489# a_13814_10483# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X57 a_293_14841# a_127_14841# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X58 a_127_3207# w_62_6889# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X59 a_6964_6922# a_6332_6922# a_6332_6922# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.32 as=0.33 ps=2.32 w=0.5 l=2.5
X60 a_12993_7763# a_12402_7915# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X61 a_12231_1209# a_12402_1387# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X62 a_13887_14265# a_14090_14543# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X63 w_62_2537# a_2371_2689# a_2539_2591# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X64 a_2073_14291# a_2038_14543# a_1835_14265# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X65 w_62_12329# a_2754_12267# a_3250_12481# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X66 a_4575_15567# a_3746_14835# a_4825_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X67 a_127_3207# div_fb2_2 a_2245_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X68 w_62_15593# a_14755_13747# a_14806_15067# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X69 a_14494_9217# a_14407_8993# a_14090_9103# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X70 a_14806_12267# a_13835_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X71 w_62_10153# a_15188_11545# a_15126_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X72 a_12353_2573# a_12265_2475# a_12271_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X73 a_397_7763# a_534_7943# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X74 a_13185_15379# a_1225_15531# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X75 a_3746_9395# a_3660_9627# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X76 a_127_3207# a_122_8539# a_127_9401# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X77 w_62_10153# a_15123_10483# a_15289_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X78 a_2313_13025# a_1835_12633# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X79 a_2442_8129# a_2355_7905# a_2038_8015# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X80 a_12586_1415# a_13435_2083# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X81 a_122_8539# a_1225_10091# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X82 a_15126_513# a_14407_289# a_14563_384# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X83 a_446_399# a_350_1387# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X84 a_14079_8281# a_13835_7763# a_14465_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X85 a_2272_14657# a_1835_14265# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X86 a_127_3207# a_6422_13265# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X87 a_774_11937# a_121_10748# a_350_11803# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X88 a_4137_292# enb_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X89 a_2245_1011# a_1783_147# a_535_2475# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X90 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=41.8133 ps=361.1 w=0.87 l=0.59
X91 w_62_7977# a_12854_9939# a_14708_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X92 a_127_3207# a_14368_9119# a_14407_8993# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X93 w_62_14505# a_2316_14559# a_2355_14433# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X94 a_127_3207# a_947_11001# a_2073_13025# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X95 a_3079_2145# a_2703_691# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X96 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X97 a_127_3207# a_11279_8265# a_11279_8265# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.225 pd=1.8 as=0.45 ps=3.6 w=1.5 l=0.15
X98 a_14873_1235# a_14494_1601# a_14801_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X99 a_127_3207# a_1383_8611# a_1317_8685# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X100 a_727_15353# a_534_14471# a_1397_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X101 a_127_3207# a_13199_8013# a_12499_10091# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X102 a_127_3207# a_947_11001# a_905_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X103 a_14365_1235# a_13887_1209# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X104 a_127_3207# a_2316_8031# a_2355_7905# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X105 w_62_9065# a_2316_9119# a_2355_8993# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X106 a_548_15201# a_127_14291# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X107 a_861_13721# a_643_14125# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X108 w_62_10153# a_15188_9100# a_15126_9217# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X109 w_62_9065# a_534_9031# a_1397_9101# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X110 a_14732_15629# a_14407_15647# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X111 w_62_14505# div_fb3_3 a_2057_14835# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X112 a_12449_13203# a_12402_13355# a_12231_13177# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X113 a_1673_10489# a_1507_10489# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X114 a_3140_1779# a_1783_1235# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X115 a_1562_11027# a_947_11001# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X116 a_11658_8851# a_11382_8851# a_11300_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X117 a_9193_4818# a_6332_5146# a_8019_5400# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.15 ps=1.3 w=1 l=0.5
X118 a_3136_13452# a_3250_13747# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X119 a_12695_12115# a_12179_12115# a_12600_12115# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X120 a_15289_9939# a_15123_9939# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X121 a_14563_384# a_14368_415# a_14873_147# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X122 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X123 a_127_3207# a_3763_11545# a_5003_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X124 w_62_7977# a_3136_8012# a_3074_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X125 a_12345_12115# a_12179_12115# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X126 a_14109_11277# a_14079_11212# a_12265_10715# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X127 a_5679_15567# a_5419_15353# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X128 w_62_361# a_122_923# a_127_697# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X129 a_14873_11937# a_14494_11571# a_14801_11937# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X130 a_127_3207# a_6422_7825# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=6
X131 a_14079_11212# a_13835_11571# a_14465_11277# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X132 w_62_361# div_fb2_0 a_2057_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X133 a_3746_1779# a_3660_2011# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X134 a_13449_147# div_out1_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X135 a_127_3207# a_121_2297# a_397_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X136 w_62_361# a_14806_923# a_15302_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X137 a_127_3207# a_6422_7825# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X138 a_12595_2297# a_12586_1415# a_13449_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X139 a_3746_14835# a_3660_15067# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X140 a_127_3207# a_7331_4818# a_12296_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X141 a_673_15629# a_631_15531# a_567_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X142 a_4533_2573# a_3899_2573# a_4315_2297# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X143 a_2038_9103# a_2355_8993# a_2313_8851# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X144 a_15302_691# a_14806_923# a_15131_1057# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X145 a_11382_11571# a_11296_11803# a_11300_11891# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X146 a_535_10715# a_2027_12300# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X147 a_13260_15213# a_12179_14841# a_12913_14809# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X148 a_127_3207# a_13835_12659# a_15131_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X149 a_12345_8313# a_12179_8313# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X150 a_127_3207# div_out0_1 a_13199_9101# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X151 a_1383_14051# a_947_14025# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X152 a_861_14809# a_643_15213# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X153 a_3763_11545# a_5003_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X154 w_62_2537# a_7331_5294# a_6332_5146# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X155 a_13887_8825# a_14090_9103# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X156 a_127_3207# a_13835_7763# a_15131_8673# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X157 a_14090_13455# a_14368_13471# a_14324_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X158 a_9567_4858# a_10437_4858# sky130_fd_pr__cap_mim_m3_1 l=6 w=7
X159 a_127_3207# a_947_969# a_2073_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X160 a_127_3207# a_179_8825# a_127_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X161 a_534_12899# a_1383_12089# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X162 w_62_10153# a_12595_9913# a_12541_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X163 a_14368_13471# a_12174_13979# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X164 w_62_7977# a_947_8585# a_2656_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X165 a_739_9773# a_127_9401# a_643_9773# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X166 w_62_10153# a_3519_10499# a_3379_10821# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X167 a_2057_8307# a_1783_7763# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X168 a_14806_923# a_13835_147# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X169 a_751_691# a_293_697# a_643_1069# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X170 a_905_8673# a_861_8281# a_739_8685# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X171 w_62_12329# a_13260_12115# a_13435_12089# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X172 a_122_11179# a_1225_10715# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X173 a_5853_11873# a_3746_12115# a_5678_11285# w_62_11241# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X174 a_534_11811# a_1383_11001# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X175 a_127_3207# a_14563_12633# a_14494_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X176 w_62_2537# a_14368_1503# a_14407_1377# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X177 a_12826_11937# a_11989_10748# a_12402_11803# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X178 w_62_7977# a_13887_7737# a_13835_7763# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X179 a_567_10189# a_535_10091# a_485_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X180 w_62_15593# a_11279_13367# a_11279_13367# w_62_15593# sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.3 as=0.9 ps=6.6 w=3 l=0.15
X181 a_127_3207# a_11989_9913# a_12449_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X182 a_127_3207# a_2114_10457# a_2072_10861# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X183 w_62_14505# a_122_13979# a_127_14841# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X184 a_127_3207# a_534_11811# a_774_11937# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X185 a_1225_2475# enb_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X186 a_127_3207# a_15123_9939# a_15289_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X187 a_127_3207# a_12854_10483# a_12957_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X188 w_62_2537# a_2114_2435# a_2041_2689# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X189 a_127_3207# a_13887_14265# a_13835_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X190 a_5225_14701# a_4971_13388# a_4971_13388# w_62_14505# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1 as=0.15 ps=1.6 w=0.5 l=0.15
X191 a_3136_1484# a_3250_1779# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X192 a_12595_9913# a_13199_9101# a_13449_9101# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X193 a_12600_15201# a_12179_14291# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X194 a_127_3207# a_1225_2475# a_5175_432# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X195 w_62_2537# a_15123_2323# a_15289_2323# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X196 w_62_14505# a_1383_15139# a_1370_14835# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X197 a_5853_13858# a_3746_13747# a_5678_14627# w_62_14505# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X198 a_1147_1485# a_534_1415# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X199 w_62_13417# div_fb1_3 a_1229_13453# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X200 a_14368_12775# a_12174_11179# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X201 a_127_3207# a_14407_2591# a_14838_2645# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X202 a_3657_9939# a_3379_9967# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X203 a_15289_10483# a_15123_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X204 a_2057_691# a_2027_665# a_535_2475# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X205 a_127_3207# a_14806_923# a_14755_691# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X206 a_14368_9119# a_12174_8539# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X207 a_14368_8031# a_12174_8539# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X208 w_62_10153# a_3519_9941# a_3379_9967# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X209 a_13369_11027# a_12345_11027# a_13260_11027# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X210 a_534_13383# a_1383_14051# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X211 a_127_3207# a_2316_13471# a_2355_13345# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X212 a_2041_2689# a_1507_2323# a_1946_2689# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X213 a_13614_1057# a_12854_2323# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X214 a_127_3207# a_4575_10457# a_4315_10457# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X215 a_4077_7948# a_4077_7948# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X216 a_12498_399# a_12402_1387# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X217 a_3136_11545# a_3250_11393# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X218 a_548_9761# a_127_8851# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X219 a_1673_9939# a_1507_9939# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X220 a_14079_14809# div_out3_3 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X221 w_62_7977# a_14563_8000# a_14494_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X222 a_1397_14291# div_fb0_3 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X223 a_127_3207# a_8169_4818# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=2
X224 a_5003_10189# a_2864_10189# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X225 w_62_2537# a_5679_2511# a_5637_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X226 a_127_3207# a_15188_13452# a_15126_13569# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X227 a_534_327# a_1383_995# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X228 a_11300_8851# a_11279_8265# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.45 pd=3.6 as=0.225 ps=1.8 w=1.5 l=0.15
X229 w_62_15593# a_14239_15745# a_14407_15647# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X230 a_13909_10483# a_13375_10489# a_13814_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X231 a_127_3207# a_403_10483# a_1507_10489# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X232 a_14090_12791# a_14368_12775# a_14324_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X233 a_2027_9369# a_1783_8851# a_2413_9395# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X234 a_4575_10127# a_4315_9913# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X235 a_127_3207# w_62_4713# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X236 a_14563_384# a_14407_289# a_14708_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X237 a_127_3207# a_12174_13979# a_12179_13753# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X238 a_127_3207# a_5853_8418# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=3.3 pd=22.6 as=0 ps=0 w=11 l=2
X239 a_127_3207# a_12174_8539# a_12179_8313# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X240 w_62_15593# a_1371_15353# a_122_13979# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X241 a_13435_9699# a_13260_9773# a_13614_9761# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X242 a_3746_12115# a_3617_11803# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X243 a_127_3207# a_122_923# a_127_1785# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X244 a_127_3207# a_7331_4818# a_8109_7110# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X245 w_62_10153# a_12595_10457# a_12541_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X246 a_5003_15629# a_2864_15629# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X247 a_121_10748# w_62_10153# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X248 a_861_8281# a_643_8685# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X249 a_4575_10457# a_4315_10457# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X250 a_3746_8307# a_3617_9003# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X251 a_2371_10483# a_1673_10489# a_2114_10457# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X252 a_397_7763# a_350_7915# a_179_7737# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X253 a_1383_8611# a_1208_8685# a_1562_8673# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X254 a_3074_1601# a_2316_1503# a_2511_1472# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X255 a_3746_11027# a_3660_11179# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X256 a_12913_9369# a_12695_9773# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X257 a_350_13355# a_446_13455# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X258 a_3136_396# a_3250_691# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X259 a_727_9913# a_1147_9101# a_1397_9101# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X260 a_13449_7763# div_out1_1 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X261 a_548_9761# a_127_8851# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X262 a_1946_10305# a_1507_9939# a_1861_9939# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X263 a_127_3207# a_14368_1503# a_14407_1377# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X264 w_62_1449# a_1225_2475# a_4971_332# w_62_1449# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1 as=0.15 ps=1.6 w=0.5 l=0.15
X265 a_5679_2511# a_5419_2297# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X266 a_567_10483# a_535_10715# a_485_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X267 a_2073_147# a_2038_399# a_1835_121# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X268 a_14090_11703# a_14368_11687# a_14324_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X269 a_127_3207# a_1383_995# a_1317_1069# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X270 a_643_8685# a_127_8313# a_548_8673# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X271 a_3899_10189# a_3657_9939# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X272 a_13909_2689# a_13375_2323# a_13814_2689# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X273 a_548_2145# a_127_1235# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X274 w_62_15593# a_15123_15379# a_15289_15379# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X275 a_127_3207# a_12586_11811# a_12826_11937# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X276 a_127_3207# a_13982_15491# a_13940_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X277 a_13260_11027# a_12345_11027# a_12913_11269# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X278 w_62_7977# a_14806_8539# a_14755_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X279 w_62_7977# a_534_7943# a_476_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X280 a_127_3207# a_1225_10715# a_5175_12724# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X281 a_12345_13753# a_12179_13753# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X282 a_15188_12633# a_15302_12481# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X283 w_62_15593# a_12913_14809# a_12803_14835# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X284 a_11658_1235# a_11382_1235# a_11300_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X285 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X286 a_548_12115# a_127_12659# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X287 a_2027_1753# a_1783_1235# a_2413_1779# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X288 a_11684_6622# a_11630_6516# a_7331_5294# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X289 a_13369_8685# a_12345_8313# a_13260_8685# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X290 w_62_9065# div_fb0_1 a_1229_9101# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X291 a_3657_10483# a_3379_10821# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X292 a_11658_11571# a_11382_11571# a_11300_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X293 w_62_2537# a_11989_2297# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X294 w_62_361# a_947_969# a_2656_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X295 a_1383_9699# a_947_8585# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X296 a_127_3207# a_2754_13979# a_2703_13747# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X297 a_14239_15745# a_13375_15379# a_13982_15491# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X298 a_5175_432# a_4971_332# a_4077_332# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X299 a_9887_6368# a_9193_6328# a_8199_7110# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.21 pd=2.21 as=0.3 ps=2.3 w=2 l=0.5
X300 a_3746_13747# a_3617_14443# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X301 a_751_8307# a_293_8313# a_643_8685# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X302 a_2027_9369# div_fb3_1 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X303 a_10073_5400# a_9567_4858# a_10437_4858# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.65 pd=2.65 as=0.6 ps=4.6 w=2 l=0.5
X304 a_534_7943# a_1383_8611# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X305 a_13422_11393# a_12179_11027# a_13260_11027# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X306 a_5853_13858# a_6422_13265# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X307 a_446_13455# a_350_14443# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X308 a_127_3207# div_out1_0 a_13199_397# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X309 a_127_3207# a_1835_8825# a_1783_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X310 w_62_14505# a_2511_14528# a_2442_14657# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X311 w_62_15593# a_12231_14265# a_12179_14291# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X312 a_15302_691# a_12993_147# a_15192_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X313 a_12826_8851# a_11989_9913# a_12402_9003# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X314 a_11296_11803# a_11658_11571# a_11300_11891# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X315 a_2038_1487# a_2355_1377# a_2313_1235# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X316 a_3250_13747# a_941_13203# a_3140_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X317 a_127_3207# a_6422_11089# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=6
X318 a_14932_15201# a_13835_14291# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X319 a_127_3207# a_6422_209# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X320 a_941_13203# a_350_13355# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X321 w_62_2537# a_7331_5294# a_7331_5294# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X322 a_127_3207# a_11296_11803# a_11903_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X323 a_15188_14540# a_15302_14835# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X324 a_127_3207# div_out0_0 a_13199_1485# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X325 a_127_3207# a_12231_13177# a_12179_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X326 a_127_3207# a_6422_7825# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=6
X327 a_1229_13453# a_534_13383# a_1147_13453# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X328 a_127_3207# a_12231_7737# a_12179_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X329 a_12586_14471# a_13435_15139# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X330 a_14563_14528# a_14368_14559# a_14873_14291# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X331 w_62_12329# a_12586_12899# a_13449_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X332 a_127_3207# a_13835_147# a_15131_1057# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X333 a_2864_2573# a_2539_2591# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X334 a_4273_10189# a_3899_10189# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X335 a_1861_9939# a_1766_10159# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X336 w_62_10153# a_727_9913# a_673_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X337 a_127_3207# div_fb1_2 a_1147_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X338 a_3660_11179# a_3763_11545# a_3709_11891# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X339 a_14465_12365# div_out2_2 w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X340 a_127_3207# a_179_1209# a_127_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X341 a_631_15531# a_1147_13453# a_1397_13453# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X342 a_14732_10189# a_14407_10207# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X343 a_4150_14088# a_4711_14627# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X344 w_62_2537# a_14239_2689# a_14407_2591# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X345 a_127_3207# a_6422_7825# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X346 a_127_3207# a_121_15353# a_397_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X347 a_739_2157# a_127_1785# a_643_2157# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X348 w_62_10153# a_15123_9939# a_15289_9939# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X349 w_62_12329# a_14806_12267# a_15302_12481# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X350 a_14125_14291# a_14090_14543# a_13887_14265# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X351 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X352 a_905_1057# a_861_665# a_739_1069# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X353 w_62_14505# a_534_14471# a_350_14443# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X354 a_350_12891# a_446_12633# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X355 a_14932_9761# a_13835_8851# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X356 a_14079_11212# div_out3_2 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X357 a_1383_2083# a_947_969# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X358 w_62_10153# a_1225_10091# a_11279_7927# w_62_10153# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X359 w_62_10153# a_403_10189# a_1507_9939# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X360 a_3079_12115# a_941_12659# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X361 a_2880_12115# a_1783_12659# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X362 a_127_3207# a_6422_11089# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X363 a_14563_9088# a_14407_8993# a_14708_9217# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X364 a_127_3207# a_11989_2297# a_12449_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X365 a_127_3207# a_1147_14541# a_727_15353# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X366 a_1861_15379# a_1766_15599# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X367 a_2749_11937# a_947_11001# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X368 a_14324_14657# a_13887_14265# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X369 w_62_10153# a_12586_11811# a_13449_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X370 a_13199_14541# a_12586_14471# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X371 w_62_14505# a_3136_14540# a_3074_14657# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X372 a_127_3207# div_fb0_2 a_1147_11571# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X373 a_14365_11937# a_13887_11545# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X374 a_11279_10695# a_5853_11873# a_11279_12307# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.225 pd=2.1 as=0.1125 ps=1.05 w=0.75 l=0.15
X375 a_127_3207# a_12854_10483# a_14125_13025# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X376 a_2511_8000# a_2355_7905# a_2656_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X377 a_4077_12724# a_1225_10715# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.125 ps=1 w=0.5 l=0.15
X378 w_62_15593# a_14368_14559# a_14407_14433# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X379 w_62_13417# a_1835_13177# a_1783_13203# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X380 a_14806_8539# a_13835_7763# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X381 w_62_9065# a_1383_9699# a_1370_9395# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X382 a_127_3207# a_3617_1387# a_3899_2573# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X383 w_62_3625# a_127_3207# w_62_3625# w_62_3625# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X384 a_9887_4858# a_9193_4818# a_8199_5400# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.105 pd=1.21 as=0.15 ps=1.3 w=1 l=0.5
X385 a_127_3207# a_14732_10189# a_15123_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X386 a_122_8539# a_1371_9913# a_1317_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X387 a_122_13979# a_1225_15531# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X388 a_12600_14113# a_12179_13203# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X389 a_4137_292# a_4137_292# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.15 ps=1.3 w=1 l=1
X390 w_62_12329# a_861_12357# a_751_12481# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X391 a_13260_12115# a_12179_12115# a_12913_12357# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X392 w_62_10153# a_14755_12115# a_14806_11179# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X393 a_350_11803# a_121_10748# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X394 w_62_2537# a_15123_2323# a_15289_2323# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X395 a_8019_4858# a_9193_4818# a_9151_5400# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.21 ps=2.21 w=2 l=0.5
X396 a_13614_11027# a_12854_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X397 a_14465_13747# div_out2_3 w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X398 a_127_3207# a_12127_10457# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X399 w_62_13417# a_534_13383# a_476_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X400 a_12993_147# a_12402_299# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X401 w_62_2537# a_7331_5294# a_6332_5146# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X402 a_3140_12481# a_1783_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X403 w_62_10153# a_2539_10457# a_2970_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X404 a_8199_7110# a_6485_6328# a_9567_6368# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=0.5
X405 a_2754_15067# a_1783_14291# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X406 a_397_11937# a_534_11811# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X407 a_12498_13455# a_12402_14443# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X408 a_12957_8673# a_12913_8281# a_12791_8685# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X409 w_62_14505# a_2703_13747# a_2754_15067# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X410 a_2316_11687# a_122_11179# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X411 a_14494_513# a_14368_415# a_14090_399# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X412 a_127_3207# a_13435_11001# a_13369_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X413 w_62_10153# a_13260_9773# a_13435_9699# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X414 a_15289_15379# a_15123_15379# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X415 a_12803_9395# a_12854_9939# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X416 a_2371_10305# a_1507_9939# a_2114_10051# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X417 w_62_11241# a_2754_11179# a_2703_11027# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X418 a_127_3207# a_3660_7915# a_5853_8418# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X419 a_2245_12115# a_1783_12659# a_535_10715# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X420 a_1397_8013# div_fb1_1 w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X421 a_2041_10305# a_1507_9939# a_1946_10305# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X422 a_12993_13203# a_12402_13355# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X423 a_127_3207# a_534_327# a_774_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X424 a_548_11027# a_127_11571# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X425 a_127_3207# a_1147_397# a_631_2475# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X426 a_127_3207# a_1783_12659# a_2027_12300# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X427 a_4273_10483# a_3899_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X428 a_4137_7908# a_4137_7908# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.15 ps=1.3 w=1 l=1
X429 w_62_10153# a_727_10457# a_673_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X430 a_127_3207# a_12174_923# a_12179_697# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X431 a_127_3207# a_1783_7763# a_2027_8281# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X432 a_643_14125# a_293_13753# a_548_14113# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X433 a_13435_2083# a_13260_2157# a_13614_2145# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X434 a_12403_10715# a_14079_12300# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X435 a_397_2475# a_2027_1753# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X436 a_5085_2573# a_2864_2573# a_5003_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X437 a_947_14025# a_403_15629# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X438 a_5419_15353# a_5003_15629# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X439 w_62_12329# a_179_12633# a_127_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X440 w_62_9065# div_fb3_1 a_2057_9395# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X441 a_3617_9003# a_4315_9913# a_4273_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X442 a_13435_14051# a_12854_15379# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X443 a_127_3207# a_14239_2689# a_14407_2591# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X444 a_13449_1485# div_out0_0 w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X445 w_62_1449# a_1383_2083# a_1370_1779# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X446 a_127_3207# a_9097_5098# a_11684_6622# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X447 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X448 w_62_10153# a_15123_10483# a_15289_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X449 a_127_3207# a_2539_15647# a_2970_15701# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X450 a_5853_8418# a_3746_8307# a_5678_9187# w_62_9065# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X451 a_127_3207# a_2371_10483# a_2539_10457# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X452 a_1383_995# a_1208_1069# a_1562_1057# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X453 a_12402_14443# a_11989_15353# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X454 a_12586_12899# a_13435_12089# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X455 w_62_9065# a_2754_9627# a_2703_9395# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X456 w_62_10153# a_14407_10207# a_14323_10305# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X457 w_62_15593# a_12586_14471# a_12402_14443# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X458 w_62_10153# a_2114_10051# a_2041_10305# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X459 a_1673_2323# a_1507_2323# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X460 a_1383_12089# a_1208_12115# a_1562_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X461 a_127_3207# a_12498_399# a_12449_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X462 a_548_2145# a_127_1235# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X463 a_13541_9939# a_13375_9939# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X464 a_1766_10159# a_2970_10261# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X465 a_2057_14835# a_1783_14291# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X466 a_2073_13025# a_2038_12791# a_1835_12633# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X467 a_12586_11811# a_13435_11001# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X468 a_2754_12267# a_941_12659# a_2880_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X469 w_62_15593# a_12595_15353# a_12541_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X470 a_14801_14291# a_12854_15379# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X471 a_13449_12659# div_out1_2 w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X472 w_62_1449# a_534_1415# a_350_1387# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X473 w_62_11241# a_179_11545# a_127_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X474 w_62_2537# a_13260_2157# a_13435_2083# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X475 a_2027_14809# a_1783_14291# a_2413_14835# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X476 a_1147_12659# a_534_12899# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X477 a_12803_1779# a_12854_2323# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X478 a_127_3207# w_62_3625# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X479 a_12913_9369# a_12695_9773# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X480 a_12854_10483# a_12271_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X481 a_3709_11891# a_3617_11803# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X482 a_12402_299# a_12498_399# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X483 a_8199_5400# a_6332_5146# a_9567_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.3 ps=2.6 w=1 l=0.5
X484 a_397_14291# a_350_14443# a_179_14265# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X485 a_15302_9395# a_14755_8307# a_15192_9395# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X486 a_15289_9939# a_15123_9939# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X487 a_2073_8851# a_2038_9103# a_1835_8825# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X488 a_13369_1069# a_12345_697# a_13260_1069# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X489 a_3981_2573# a_3657_2323# a_3899_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X490 a_127_3207# a_14806_12267# a_14755_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X491 a_11654_6816# a_11654_6816# a_11594_6922# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=2.1
X492 w_62_12329# a_534_12899# a_476_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X493 a_11382_1235# a_11296_1387# a_11300_1485# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X494 a_12913_665# a_12695_1069# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X495 a_567_15629# a_535_15531# a_485_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X496 w_62_15593# a_2539_15647# a_2455_15745# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X497 a_12957_15201# a_12913_14809# a_12791_15213# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X498 w_62_15593# a_13435_15139# a_13422_14835# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X499 a_2656_1601# a_2442_1601# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X500 a_127_3207# w_62_4713# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X501 a_127_3207# a_3660_12891# a_11296_11803# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X502 w_62_1449# div_fb3_0 a_2057_1779# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X503 a_127_3207# a_1783_13203# a_3079_14113# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X504 a_12271_15629# a_12265_15531# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
X505 a_127_3207# a_1835_1209# a_1783_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X506 a_941_7763# a_350_7915# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X507 a_12449_11937# a_12586_11811# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X508 a_13199_397# a_12586_327# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X509 a_12449_7763# a_12402_7915# a_12231_7737# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X510 w_62_2537# a_12231_1209# a_12179_1235# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X511 a_12826_1235# a_11989_2297# a_12402_1387# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X512 w_62_4713# a_127_3207# w_62_4713# w_62_4713# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=3.6192 ps=36.16 w=0.87 l=4.73
X513 a_12586_13383# a_13435_14051# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X514 a_13449_11571# div_out0_2 w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X515 w_62_1449# a_2754_2011# a_2703_1779# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X516 a_13260_9773# a_12345_9401# a_12913_9369# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X517 w_62_15593# a_12174_13979# a_12179_14841# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X518 a_127_3207# a_14368_13471# a_14407_13345# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X519 a_3657_15379# a_3379_15407# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X520 a_1147_11571# a_534_11811# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X521 a_3657_9939# a_3379_9967# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X522 a_861_8281# a_643_8685# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X523 a_293_14841# a_127_14841# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X524 a_15302_12481# a_14806_12267# a_15131_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X525 a_12541_10189# a_12499_10091# a_12435_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X526 a_1766_10159# a_2970_10261# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X527 w_62_15593# a_3519_15381# a_3379_15407# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X528 a_127_3207# a_1835_12633# a_1783_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X529 a_14494_8129# a_14368_8031# a_14090_8015# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X530 w_62_11241# a_534_11811# a_476_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X531 a_127_3207# a_12403_15531# a_12271_15629# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X532 w_62_5801# a_127_3207# w_62_5801# w_62_5801# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=3.6192 ps=36.16 w=0.87 l=4.73
X533 w_62_9065# a_861_9369# a_751_9395# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X534 a_12600_11027# a_12179_11571# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X535 w_62_4713# a_127_3207# w_62_4713# w_62_4713# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X536 w_62_15593# a_14806_15067# a_14755_14835# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X537 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X538 a_3709_8851# a_3617_9003# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X539 w_62_11241# a_1383_11001# a_1370_11393# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X540 a_12695_14125# a_12345_13753# a_12600_14113# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X541 a_15192_8307# a_13835_7763# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X542 a_2027_665# div_fb2_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X543 w_62_2537# a_7331_5294# a_6332_6922# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X544 w_62_7977# a_12586_7943# a_12528_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X545 a_774_14291# a_121_15353# a_350_14443# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X546 a_12913_1753# a_12695_2157# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X547 a_3617_11803# a_4315_10457# a_4273_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X548 a_127_3207# a_947_8585# a_905_8673# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X549 a_751_12481# a_947_11001# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X550 w_62_10153# a_12586_9031# a_12402_9003# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X551 a_13982_15491# a_13814_15745# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X552 a_15302_1779# a_14755_691# a_15192_1779# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X553 w_62_6889# a_127_3207# w_62_6889# w_62_6889# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=3.6192 ps=36.16 w=0.87 l=4.73
X554 a_15126_8129# a_14368_8031# a_14563_8000# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X555 a_14932_2145# a_13835_1235# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X556 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X557 a_2754_9627# a_1783_8851# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X558 w_62_361# a_12854_2323# a_14708_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X559 a_127_3207# a_14563_9088# a_14494_9217# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X560 a_1208_8685# a_293_8313# a_861_8281# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X561 a_2511_13440# a_2355_13345# a_2656_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X562 a_751_12481# a_293_12115# a_643_12115# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X563 a_2057_12365# a_2027_12300# a_535_10715# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X564 a_14109_691# a_14079_665# a_12403_2475# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X565 w_62_15593# a_11989_15353# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X566 a_13541_2323# a_13375_2323# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X567 a_2497_10861# a_1507_10489# a_2371_10483# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X568 a_127_3207# a_403_10189# a_1507_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X569 a_1766_10647# a_2970_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X570 w_62_7977# a_12586_7943# a_13449_8013# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X571 a_127_3207# a_1835_11545# a_1783_11571# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X572 a_2442_14657# a_2316_14559# a_2038_14543# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X573 a_2821_7763# a_2442_8129# a_2749_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X574 a_2272_1601# a_1835_1209# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X575 a_13260_2157# a_12345_1785# a_12913_1753# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X576 a_12803_12481# a_12854_10483# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X577 a_12402_1387# a_11989_2297# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X578 w_62_10153# a_5679_10127# a_5637_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X579 a_14873_14291# a_14494_14657# a_14801_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X580 a_2313_7763# a_1835_7737# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X581 a_14563_8000# a_14368_8031# a_14873_7763# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X582 a_14465_9395# div_out3_1 w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X583 a_127_3207# a_12595_2297# a_12271_2573# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X584 a_127_3207# a_7331_4818# a_7331_4818# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X585 w_62_13417# a_534_13383# a_1397_13453# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X586 a_11300_14541# a_11279_13367# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8 ad=0.9 pd=6.6 as=0.45 ps=3.3 w=3 l=0.15
X587 w_62_361# a_11296_1387# a_11903_147# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X588 a_12174_13979# a_1371_15353# a_13185_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X589 a_127_3207# a_3660_7915# a_11296_9003# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X590 a_15188_9100# a_15302_9395# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X591 a_127_3207# div_out2_2 a_14297_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X592 w_62_2537# a_2539_2591# a_2455_2689# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X593 a_1208_9773# a_127_9401# a_861_9369# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X594 a_15289_10483# a_15123_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X595 a_127_3207# a_13835_1235# a_14079_1753# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X596 a_2114_2435# a_1946_2689# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X597 a_4315_10457# a_3899_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X598 a_12913_12357# a_12695_12115# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X599 a_127_3207# w_62_3625# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X600 w_62_1449# a_861_1753# a_751_1779# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X601 a_2114_2435# a_1946_2689# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X602 a_5377_2573# a_5003_2573# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X603 a_6185_3321# a_9567_6368# a_10073_7110# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.325 ps=1.65 w=1 l=0.5
X604 a_548_1057# a_127_147# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X605 w_62_3625# a_127_3207# w_62_3625# w_62_3625# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X606 a_2038_14543# a_2316_14559# a_2272_14657# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X607 w_62_361# a_534_327# a_476_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X608 w_62_2537# a_14732_2573# a_15123_2323# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X609 w_62_2537# a_1371_2297# a_122_923# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X610 a_13729_9939# a_13634_10159# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X611 a_2038_9103# a_2316_9119# a_2272_9217# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X612 a_3074_513# a_2316_415# a_2511_384# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X613 a_12957_1057# a_12913_665# a_12791_1069# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X614 a_1946_15745# a_1673_15379# a_1861_15379# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X615 a_2754_2011# a_1783_1235# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X616 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X617 a_631_10091# a_534_7943# a_1397_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X618 a_127_3207# a_7331_4818# a_6485_5594# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X619 a_2057_13747# a_2027_13721# a_535_15531# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X620 w_62_15593# a_14563_14528# a_14494_14657# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X621 a_15126_14657# a_14407_14433# a_14563_14528# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X622 a_2413_8307# div_fb2_1 w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X623 a_2114_15491# a_1946_15745# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X624 a_127_3207# a_3136_11545# a_3074_11571# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X625 a_10097_3881# a_8169_4818# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X626 a_13814_15745# a_13541_15379# a_13729_15379# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X627 a_12541_10483# a_12499_10715# a_12435_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X628 a_1946_15745# a_1507_15379# a_1861_15379# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X629 a_127_3207# a_14732_10483# a_15123_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X630 w_62_15593# div_out3_3 a_14109_14835# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X631 a_15302_13747# a_12993_13203# a_15192_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X632 a_1229_8013# a_534_7943# a_1147_8013# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X633 a_14125_147# a_14090_399# a_13887_121# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X634 a_127_3207# a_1383_14051# a_1317_14125# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X635 a_127_3207# a_947_969# a_2073_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X636 a_1225_10091# a_3660_7915# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X637 w_62_10153# a_12913_11269# a_12803_11393# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X638 a_14465_1779# div_out3_0 w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X639 a_13281_9101# a_12586_9031# a_13199_9101# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X640 a_12826_14291# a_11989_15353# a_12402_14443# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X641 a_2821_13203# a_2442_13569# a_2749_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X642 a_127_3207# div_fb2_1 a_2245_8627# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X643 a_293_9401# a_127_9401# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X644 a_1208_14125# a_293_13753# a_861_13721# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X645 a_4711_9187# a_4077_7948# a_4137_7908# w_62_9065# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=1
X646 a_127_3207# a_534_14471# a_774_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X647 a_2511_12633# a_2355_12901# a_2656_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X648 a_14806_8539# a_12993_7763# a_14932_8673# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X649 a_127_3207# div_out3_1 a_14297_9715# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X650 a_861_11269# a_643_11027# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X651 w_62_1449# a_947_969# a_1835_1209# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X652 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X653 a_3250_13747# a_2754_13979# a_3079_14113# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X654 a_12803_12481# a_12345_12115# a_12695_12115# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X655 w_62_361# a_534_327# a_1397_397# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X656 w_62_361# a_2511_384# a_2442_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X657 a_127_3207# a_2754_8539# a_2703_8307# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X658 a_4273_15629# a_3899_15629# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X659 w_62_2537# a_403_2573# a_1507_2323# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X660 w_62_15593# a_727_15353# a_673_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X661 a_2038_14543# a_2355_14433# a_2313_14291# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X662 a_14079_665# a_13835_147# a_14465_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X663 a_127_3207# a_122_13979# a_127_14841# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X664 a_13541_10489# a_13375_10489# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X665 a_15131_12115# a_12993_12659# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X666 w_62_361# a_14806_923# a_14755_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X667 a_5853_802# a_6422_209# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X668 w_62_15593# a_15123_15379# a_15289_15379# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X669 a_12528_513# a_12498_399# a_12231_121# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X670 w_62_13417# a_1208_14125# a_1383_14051# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X671 a_127_3207# a_5419_10457# a_3763_11545# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X672 w_62_2537# a_13238_4858# a_13835_5043# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X673 a_127_3207# a_13199_14541# a_12595_15353# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X674 w_62_10153# a_5679_10457# a_5637_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X675 a_476_1601# a_121_2297# a_179_1209# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X676 a_643_8685# a_293_8313# a_548_8673# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X677 a_2245_2099# a_1783_1235# a_397_2475# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X678 w_62_2537# a_7331_5294# a_8109_5400# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X679 a_13982_10457# a_13814_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X680 a_12913_14809# a_12695_15213# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X681 w_62_15593# a_15188_14540# a_15126_14657# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X682 a_2073_1235# a_2038_1487# a_1835_1209# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X683 a_127_3207# a_179_121# a_127_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X684 a_3074_13569# a_2355_13345# a_2511_13440# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X685 a_2511_11545# a_2355_11813# a_2656_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X686 w_62_13417# a_13887_13177# a_13835_13203# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X687 a_12174_8539# a_1371_9913# a_13185_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X688 a_3250_8307# a_2754_8539# a_3079_8673# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X689 a_2057_9395# a_2027_9369# a_397_10091# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X690 a_14090_1487# a_14368_1503# a_14324_1601# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X691 a_13238_4858# a_12183_5294# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=0.5
X692 a_643_11027# a_293_11027# a_548_11027# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X693 w_62_10153# a_11279_10695# a_11279_10695# w_62_10153# sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.3 as=0.9 ps=6.6 w=3 l=0.15
X694 a_403_10189# a_631_10091# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X695 a_4137_12618# a_3660_12891# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X696 a_127_3207# w_62_3625# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X697 a_15302_9395# a_14806_9627# a_15131_9761# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X698 a_127_3207# a_12586_9031# a_12826_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X699 a_127_3207# a_14407_10457# a_14365_10861# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X700 a_2511_13440# a_2316_13471# a_2821_13203# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X701 a_127_3207# a_6422_11089# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=6
X702 a_3899_10483# a_3657_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X703 a_6964_4858# a_6332_5146# a_6332_5146# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.32 as=0.33 ps=2.32 w=0.5 l=2.5
X704 a_10073_6368# a_9567_6368# a_6185_3321# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.65 pd=2.65 as=0.6 ps=4.6 w=2 l=0.5
X705 a_12271_10189# a_12499_10091# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X706 a_11382_14291# a_11296_14443# a_11300_14541# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X707 w_62_2537# a_12174_923# a_12179_1785# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X708 a_15192_12481# a_13835_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X709 a_259_2517# a_127_3207# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X710 a_13369_15213# a_12345_14841# a_13260_15213# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X711 a_4150_12042# a_4711_11285# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X712 a_485_10189# a_397_10091# a_403_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X713 a_1397_13453# div_fb1_3 w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X714 a_2656_13569# a_2442_13569# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X715 w_62_10153# a_14407_10457# a_14838_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X716 a_14297_12115# a_13835_12659# a_12403_10715# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X717 a_12127_2517# a_127_3207# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X718 a_631_10715# a_534_12899# a_1397_12979# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X719 a_3709_1235# a_3617_1387# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X720 a_12595_15353# a_13199_14541# a_13449_14541# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X721 w_62_361# a_1835_121# a_1783_147# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X722 a_3657_2323# a_3379_2351# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.475 pd=2.95 as=0.16655 ps=1.39 w=1 l=0.15
X723 a_127_3207# a_13238_4858# a_13835_5043# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X724 a_127_3207# a_947_969# a_905_1057# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X725 w_62_2537# clk_ref_0 a_3379_2351# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.16655 pd=1.39 as=0.0567 ps=0.69 w=0.42 l=0.15
X726 w_62_9065# a_4077_7948# a_5678_9187# w_62_9065# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X727 a_905_12115# a_861_12357# a_739_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X728 a_127_3207# a_6422_11089# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X729 a_1766_2543# a_2970_2645# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X730 a_2656_513# a_2442_513# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X731 a_127_3207# a_4137_292# a_4077_332# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.3 ps=2.6 w=1 l=1
X732 a_12528_9217# a_11989_9913# a_12231_8825# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X733 a_127_3207# a_12586_14471# a_12826_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X734 a_2057_1779# a_2027_1753# a_397_2475# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X735 w_62_7977# a_2754_8539# a_3250_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X736 a_1835_13177# a_2038_13455# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X737 a_127_3207# a_14563_1472# a_14494_1601# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X738 w_62_2537# a_11749_5294# a_11648_4958# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=0.5
X739 a_12403_10091# a_14079_8281# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X740 a_4137_292# a_4077_332# a_4711_1571# w_62_1449# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=1
X741 a_15126_9217# a_14407_8993# a_14563_9088# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X742 w_62_4713# a_127_3207# w_62_4713# w_62_4713# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X743 a_127_3207# a_13835_14291# a_14079_14809# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X744 a_2754_11179# a_1783_11571# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X745 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X746 w_62_11241# a_2703_12115# a_2754_11179# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X747 a_127_3207# w_62_5801# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X748 a_127_3207# a_3136_8012# a_3074_8129# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X749 a_3617_14443# a_4315_15353# a_4273_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X750 a_13435_12089# a_13260_12115# a_13614_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X751 a_12449_147# a_12402_299# a_12231_121# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X752 a_127_3207# a_5419_9913# a_3763_8825# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X753 a_179_13177# a_350_13355# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X754 a_1370_12481# a_127_12115# a_1208_12115# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X755 a_727_10457# a_534_11811# a_1397_11891# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X756 a_127_3207# a_14407_15647# a_14838_15701# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X757 a_2316_11687# a_122_11179# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X758 a_12913_665# a_12695_1069# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X759 a_8109_7110# a_6185_3321# a_8019_7110# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.3 ps=2.6 w=1 l=0.15
X760 w_62_7977# div_out1_1 a_13281_8013# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X761 a_1370_8307# a_127_8313# a_1208_8685# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X762 a_127_3207# a_446_12633# a_397_13025# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X763 a_14109_14835# a_13835_14291# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X764 a_941_12659# a_350_12891# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X765 a_12345_13753# a_12179_13753# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X766 a_13238_4858# a_11648_4958# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
X767 a_2442_13569# a_2355_13345# a_2038_13455# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X768 a_14125_13025# a_14090_12791# a_13887_12633# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X769 a_127_3207# a_15188_9100# a_15126_9217# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X770 a_14806_12267# a_12993_12659# a_14932_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X771 w_62_10153# a_13982_10051# a_13909_10305# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X772 w_62_12329# a_12231_12633# a_12179_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X773 a_350_9003# a_121_9913# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X774 w_62_7977# a_179_7737# a_127_7763# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X775 a_127_3207# w_62_6889# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X776 a_13614_9761# a_12854_9939# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X777 a_1208_2157# a_127_1785# a_861_1753# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X778 a_13634_10159# a_14838_10261# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X779 a_127_3207# a_3763_14265# a_5003_15629# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X780 a_14079_8281# div_out2_1 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X781 a_127_3207# a_535_2475# a_403_2573# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X782 a_1766_15599# a_2970_15701# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X783 a_127_3207# a_3746_11027# a_4575_10457# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X784 a_10073_4858# a_9567_4858# a_10437_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.325 pd=1.65 as=0.3 ps=2.6 w=1 l=0.5
X785 a_14708_8129# a_14494_8129# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X786 a_14109_9395# a_13835_8851# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X787 a_3465_9967# a_1225_10091# a_3379_9967# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X788 w_62_10153# a_12913_9369# a_12803_9395# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X789 a_13185_2323# a_1225_2475# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X790 a_12695_11027# a_12345_11027# a_12600_11027# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X791 a_1562_8673# a_947_8585# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X792 w_62_11241# a_2316_11687# a_2355_11813# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X793 a_127_3207# a_2511_384# a_2442_513# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X794 a_127_3207# a_11296_1387# a_11903_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X795 w_62_1449# a_534_1415# a_1397_1485# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X796 a_127_3207# a_13199_397# a_12499_2475# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X797 a_127_3207# a_8169_4818# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X798 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X799 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X800 a_8019_7110# a_9193_6328# a_9151_6368# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.21 ps=2.21 w=2 l=0.5
X801 a_12498_8015# a_12402_9003# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X802 a_127_3207# a_12403_2475# a_12271_2573# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X803 w_62_2537# a_7331_5294# a_6332_6922# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X804 a_13435_8611# a_12854_9939# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X805 a_127_3207# a_13835_13203# a_15131_14113# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X806 w_62_10153# a_12271_10483# a_13375_10489# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X807 a_127_3207# a_14806_2011# a_14755_1779# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X808 a_15289_15379# a_15123_15379# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X809 w_62_2537# a_2539_2591# a_2970_2645# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X810 a_643_14125# a_127_13753# a_548_14113# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X811 a_446_12633# a_350_11803# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X812 a_397_8851# a_534_9031# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X813 a_3074_13569# a_2316_13471# a_2511_13440# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X814 a_403_2573# a_397_2475# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
X815 w_62_361# a_941_147# a_2754_923# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X816 w_62_10153# a_12231_11545# a_12179_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X817 a_2656_12659# a_2442_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X818 a_15188_396# a_15302_691# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X819 a_485_10483# a_397_10715# a_403_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X820 a_2442_9217# a_2355_8993# a_2038_9103# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X821 a_14932_11027# a_13835_11571# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X822 a_12791_14125# a_12179_13753# a_12695_14125# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X823 a_5175_8048# a_4971_7948# a_4077_7948# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X824 a_127_3207# div_fb1_1 a_1147_8013# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X825 a_3763_14265# a_5003_15629# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X826 w_62_2537# a_3763_1209# a_5085_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X827 a_12271_2573# a_12265_2475# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
X828 a_1835_7737# a_2038_8015# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X829 a_11279_13705# a_3660_13355# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X830 a_3074_12659# a_2355_12901# a_2511_12633# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X831 a_2114_10457# a_1946_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X832 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X833 a_127_3207# a_13887_12633# a_13835_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X834 a_534_1415# a_1383_2083# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X835 a_3617_9003# a_3899_10189# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X836 a_14239_10483# a_13375_10489# a_13982_10457# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X837 w_62_10153# a_12854_9939# a_14708_9217# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X838 w_62_9065# a_3763_8825# a_3660_9627# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X839 w_62_3625# a_127_3207# w_62_3625# w_62_3625# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X840 a_1835_12633# a_2038_12791# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X841 a_127_3207# a_1383_9699# a_1317_9773# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X842 a_2749_14291# a_947_14025# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X843 w_62_10153# a_13435_11001# a_13422_11393# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X844 w_62_2537# a_6185_3209# a_13743_5587# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X845 a_127_3207# a_13199_9101# a_12595_9913# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X846 a_127_3207# a_947_11001# a_905_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X847 a_14365_14291# a_13887_14265# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X848 a_14109_1779# a_13835_1235# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X849 a_861_14809# a_643_15213# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X850 a_2316_415# a_122_923# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X851 w_62_2537# a_12913_1753# a_12803_1779# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X852 a_14806_923# a_12993_147# a_14932_1057# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X853 a_127_3207# a_2316_9119# a_2355_8993# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X854 a_2511_12633# a_2316_12775# a_2821_13025# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X855 a_12541_15629# a_12499_15531# a_12435_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X856 a_179_7737# a_350_7915# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X857 a_2656_11571# a_2442_11571# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X858 a_127_3207# a_1147_8013# a_631_10091# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X859 a_1562_12115# a_947_11001# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X860 w_62_13417# a_2754_13979# a_3250_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X861 a_3136_14540# a_3250_14835# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X862 a_179_12633# a_350_12891# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X863 a_14563_13440# a_14407_13345# a_14708_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X864 w_62_9065# a_3136_9100# a_3074_9217# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X865 a_14806_13979# a_13835_13203# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X866 a_127_3207# a_14563_13440# a_14494_13569# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X867 a_14465_691# div_out2_0 w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X868 a_14324_8129# a_13887_7737# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X869 a_14109_12365# a_14079_12300# a_12403_10715# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X870 a_127_3207# a_3746_9395# a_5679_10127# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X871 a_2442_12659# a_2355_12901# a_2038_12791# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X872 a_14563_11545# a_14368_11687# a_14873_11937# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X873 a_403_10483# a_631_10715# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X874 a_3763_1209# a_5003_2573# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X875 a_4971_7948# a_4137_7908# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X876 a_1397_12979# div_fb1_2 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X877 a_643_1069# a_293_697# a_548_1057# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X878 a_14079_12300# a_13835_12659# a_14465_12365# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X879 a_127_3207# a_13887_11545# a_13835_11571# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X880 a_13281_13453# a_12586_13383# a_13199_13453# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X881 a_12993_12659# a_12402_12891# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X882 a_8019_5400# a_9193_4818# a_9151_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.105 ps=1.21 w=1 l=0.5
X883 a_11300_1235# a_11279_649# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.45 pd=3.6 as=0.225 ps=1.8 w=1.5 l=0.15
X884 w_62_13417# a_12854_15379# a_14708_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X885 a_13814_2689# a_13541_2323# a_13729_2323# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X886 a_397_14291# a_534_14471# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X887 a_127_3207# a_2511_11545# a_2442_11571# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X888 a_1835_11545# a_2038_11703# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X889 a_1861_15379# a_1766_15599# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X890 a_127_3207# a_7331_4818# a_6485_5594# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X891 a_293_8313# a_127_8313# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X892 a_13634_10647# a_14838_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X893 a_14365_15379# a_13375_15379# a_14239_15745# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X894 a_3250_691# a_2754_923# a_3079_1057# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X895 w_62_10153# a_11279_7927# a_11279_7927# w_62_10153# sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.3 as=0.9 ps=6.6 w=3 l=0.15
X896 a_2072_15379# a_1673_15379# a_1946_15745# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X897 a_127_3207# div_out2_0 a_14297_1011# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X898 a_127_3207# a_11989_10748# a_12449_11937# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X899 w_62_7977# a_13435_8611# a_13422_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X900 a_4150_12042# a_4910_12154# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X901 a_2316_8031# a_122_8539# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X902 a_127_3207# a_13835_11571# a_14079_11212# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X903 a_15302_1779# a_14806_2011# a_15131_2145# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X904 a_12595_2297# a_13199_1485# a_13449_1485# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X905 a_13982_2435# a_13814_2689# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X906 a_12435_10189# a_12403_10091# a_12353_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X907 a_127_3207# a_4575_15567# a_4315_15353# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X908 a_127_3207# a_12586_1415# a_12826_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X909 a_179_11545# a_350_11803# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X910 a_12345_9401# a_12179_9401# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X911 a_11296_14443# a_11658_14291# a_11300_14541# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X912 a_14801_13025# a_12854_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X913 w_62_15593# a_5679_15567# a_5637_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X914 a_774_147# a_446_399# a_350_299# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X915 a_15188_8012# a_15302_8307# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X916 a_1383_15139# a_947_14025# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X917 a_5679_10127# a_3746_9395# a_5929_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X918 w_62_2537# a_1371_2297# a_12174_923# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X919 a_14494_1601# a_14407_1377# a_14090_1487# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X920 a_127_3207# a_13835_8851# a_15131_9761# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X921 a_3074_12659# a_2316_12775# a_2511_12633# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X922 a_2442_11571# a_2355_11813# a_2038_11703# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X923 a_14090_14543# a_14368_14559# a_14324_14657# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X924 a_127_3207# a_4137_13348# a_4077_13388# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.3 ps=2.6 w=1 l=1
X925 a_127_3207# div_out0_3 a_13199_14541# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X926 a_4315_2297# a_3899_2573# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X927 a_673_2573# a_631_2475# a_567_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X928 a_13743_5587# a_6185_3209# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X929 a_2313_13203# a_1835_13177# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X930 a_1397_11891# div_fb0_2 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X931 a_12296_4858# a_7331_4818# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X932 a_12498_12633# a_12402_11803# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X933 a_14368_14559# a_12174_13979# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X934 a_12695_14125# a_12179_13753# a_12600_14113# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X935 w_62_9065# a_947_8585# a_2656_9217# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X936 a_397_13025# a_350_12891# a_179_12633# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X937 a_127_3207# a_1783_7763# a_3079_8673# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X938 a_259_10133# a_127_3207# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X939 w_62_14505# a_3763_14265# a_3660_15067# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X940 a_293_11027# a_127_11027# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X941 a_8199_7110# a_5853_802# a_8109_7110# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.15 ps=1.3 w=1 l=0.15
X942 a_905_9761# a_861_9369# a_739_9773# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X943 a_12541_2573# a_12499_2475# a_12435_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X944 a_14365_2323# a_13375_2323# a_14239_2689# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X945 a_14109_13747# a_14079_13721# a_12403_15531# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X946 a_127_3207# a_947_14025# a_2073_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X947 a_534_12899# a_1383_12089# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X948 a_2027_13721# div_fb2_3 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X949 a_2864_2573# a_2539_2591# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X950 a_14079_13721# a_13835_13203# a_14465_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X951 a_127_3207# a_3617_11803# a_3899_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X952 a_127_3207# w_62_3625# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X953 w_62_10153# a_13887_8825# a_13835_8851# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X954 a_4575_15567# a_4315_15353# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X955 w_62_361# a_534_327# a_350_299# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X956 w_62_2537# a_7331_5294# a_8109_5400# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X957 a_12586_9031# a_13435_9699# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X958 a_3074_11571# a_2316_11687# a_2511_11545# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X959 a_127_3207# a_12854_10483# a_12957_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X960 a_2316_415# a_122_923# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X961 a_127_3207# a_14407_2591# a_14365_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X962 w_62_1449# a_2316_1503# a_2355_1377# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X963 w_62_7977# a_12854_9939# a_13887_7737# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X964 w_62_2537# a_13982_2435# a_13909_2689# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X965 a_15126_1601# a_14407_1377# a_14563_1472# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X966 w_62_7977# a_1835_7737# a_1783_7763# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X967 w_62_2537# a_15188_1484# a_15126_1601# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X968 a_6185_3881# a_9585_3657# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X969 w_62_3625# a_127_3207# w_62_3625# w_62_3625# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X970 w_62_14505# div_fb0_3 a_1229_14541# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X971 a_14563_12633# a_14407_12901# a_14708_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X972 a_2455_10305# a_1673_9939# a_2371_10305# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X973 a_4825_2573# a_4315_2297# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X974 a_548_14113# a_127_13203# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X975 a_1397_397# div_fb1_0 w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X976 a_14368_9119# a_12174_8539# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X977 w_62_12329# a_12854_10483# a_14708_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X978 a_127_3207# a_2539_15647# a_2497_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X979 a_774_13025# a_446_12633# a_350_12891# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X980 a_127_3207# a_15123_2323# a_15289_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X981 a_15126_513# a_14368_415# a_14563_384# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X982 w_62_7977# div_out2_1 a_14109_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X983 a_127_3207# div_fb1_3 a_1147_13453# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X984 a_13369_12115# a_12345_12115# a_13260_12115# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X985 a_127_3207# a_15188_1484# a_15126_1601# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X986 a_727_2297# a_1147_1485# a_1397_1485# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X987 a_14323_10305# a_13541_9939# a_14239_10305# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X988 a_534_14471# a_1383_15139# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X989 a_5175_13488# a_4971_13388# a_4077_13388# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X990 a_127_3207# a_1225_10091# a_5175_8048# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X991 a_3617_11803# a_3899_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X992 a_13614_2145# a_12854_2323# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X993 w_62_13417# a_13260_14125# a_13435_14051# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X994 a_3136_12633# a_3250_12481# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X995 a_12449_14291# a_12586_14471# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X996 a_12449_7763# a_12586_7943# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X997 w_62_7977# a_122_8539# a_127_8313# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X998 a_3763_1209# a_5419_2297# a_5377_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X999 a_2864_10483# a_2539_10457# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1000 a_10073_7110# a_9097_5098# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.325 ps=1.65 w=1 l=0.15
X1001 w_62_10153# a_14563_9088# a_14494_9217# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1002 a_122_11179# a_1371_10457# a_1317_10803# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1003 a_4150_8648# a_4711_9187# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X1004 a_12957_11027# a_12913_11269# a_12791_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1005 a_397_147# a_534_327# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1006 a_1562_1057# a_947_969# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1007 a_14297_8627# a_13835_7763# a_12403_10091# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X1008 a_14563_11545# a_14407_11813# a_14708_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1009 a_12174_8539# a_1225_10091# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1010 a_127_3207# a_11279_649# a_11279_649# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.225 pd=1.8 as=0.45 ps=3.6 w=1.5 l=0.15
X1011 w_62_10153# a_2371_10305# a_2539_10207# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1012 a_3136_11545# a_3250_11393# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1013 a_12498_399# a_12402_1387# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1014 a_12435_10483# a_12403_10715# a_12353_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X1015 a_2821_147# a_2442_513# a_2749_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1016 a_127_3207# a_12854_2323# a_14125_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1017 w_62_7977# a_2511_8000# a_2442_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1018 w_62_1449# div_fb0_0 a_1229_1485# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1019 a_5679_10457# a_3746_11027# a_5929_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1020 a_13887_1209# a_14090_1487# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1021 a_127_3207# w_62_5801# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1022 a_12586_1415# a_13435_2083# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1023 a_127_3207# a_12174_13979# a_12179_14841# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1024 a_14873_13025# a_14494_12659# a_14801_13025# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1025 w_62_10153# a_12854_10483# a_14708_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1026 a_127_3207# a_12174_8539# a_12179_9401# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1027 a_2057_691# a_1783_147# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1028 a_397_1235# a_534_1415# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1029 a_1225_15531# a_3660_13355# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1030 a_6185_3209# a_9585_3209# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X1031 a_4150_1032# a_4910_920# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X1032 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1033 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1034 a_861_9369# a_643_9773# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1035 a_12791_8685# a_12179_8313# a_12695_8685# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1036 a_293_11027# a_127_11027# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1037 a_3746_9395# a_3660_9627# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1038 a_127_3207# a_1147_12659# a_631_10715# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1039 w_62_361# a_14563_384# a_14494_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1040 a_397_8851# a_350_9003# a_179_8825# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1041 a_1383_9699# a_1208_9773# a_1562_9761# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1042 a_2371_10305# a_1673_9939# a_2114_10051# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1043 a_127_3207# a_15123_10483# a_15289_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1044 a_13541_10489# a_13375_10489# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1045 a_13199_12659# a_12586_12899# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1046 a_12803_691# a_12854_2323# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1047 a_127_3207# enb_0 a_7331_4818# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X1048 a_3746_12115# a_3617_11803# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1049 w_62_10153# a_2539_10457# a_2455_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1050 a_350_14443# a_121_15353# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X1051 a_13449_8851# div_out0_1 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1052 a_12449_11937# a_12402_11803# a_12231_11545# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1053 a_14708_13569# a_14494_13569# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1054 a_3079_14113# a_941_13203# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1055 a_15131_8673# a_12993_7763# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1056 a_11300_9101# a_11279_7927# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8 ad=0.9 pd=6.6 as=0.45 ps=3.3 w=3 l=0.15
X1057 a_127_3207# a_1383_2083# a_1317_2157# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1058 a_2880_14113# a_1783_13203# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X1059 a_127_3207# a_13199_1485# a_12595_2297# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1060 a_3136_13452# a_3250_13747# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X1061 a_485_15629# a_397_15531# a_403_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X1062 a_127_3207# a_2316_1503# a_2355_1377# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1063 a_4077_7948# a_1225_10091# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.125 ps=1 w=0.5 l=0.15
X1064 a_11989_10748# w_62_10153# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1065 a_4971_332# a_4137_292# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X1066 w_62_2537# a_14563_1472# a_14494_1601# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1067 a_2880_8673# a_1783_7763# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X1068 a_13260_12115# a_12345_12115# a_12913_12357# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1069 w_62_9065# a_534_9031# a_476_9217# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X1070 a_12345_14841# a_12179_14841# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1071 a_14368_13471# a_12174_13979# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1072 a_2413_11277# div_fb3_2 w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1073 w_62_2537# a_6185_3209# a_13743_5587# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1074 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1075 a_127_3207# a_2511_14528# a_2442_14657# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1076 a_127_3207# a_1147_11571# a_727_10457# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1077 a_13369_9773# a_12345_9401# a_13260_9773# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1078 a_3660_15067# a_3617_14443# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1079 a_13199_11571# a_12586_11811# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1080 a_4077_13388# a_1225_15531# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.125 ps=1 w=0.5 l=0.15
X1081 w_62_12329# a_4910_12154# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X1082 w_62_11241# a_122_11179# a_127_11027# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1083 w_62_361# div_out2_0 a_14109_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1084 a_13729_15379# a_13634_15599# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1085 a_14368_1503# a_12174_923# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1086 a_127_3207# a_2754_15067# a_2703_14835# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1087 a_127_3207# a_6422_209# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X1088 a_12826_13025# a_12498_12633# a_12402_12891# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1089 a_3746_14835# a_3660_15067# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1090 w_62_361# a_12993_147# a_14806_923# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X1091 a_3136_9100# a_3250_9395# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X1092 a_127_3207# div_fb2_3 a_2245_14067# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1093 a_15289_9939# a_15123_9939# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1094 a_13422_12481# a_12179_12115# a_13260_12115# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1095 a_4077_332# a_4077_332# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X1096 a_127_3207# a_534_12899# a_774_13025# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X1097 a_293_697# a_127_697# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1098 a_12791_11027# a_12179_11027# a_12695_11027# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1099 a_127_3207# a_11654_6816# a_12074_7210# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X1100 w_62_2537# a_7331_5294# a_8109_6368# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X1101 a_11382_8851# a_11296_9003# a_11300_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1102 a_5853_8418# a_3763_8825# a_5678_8030# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X1103 a_127_3207# a_4137_292# a_5678_414# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X1104 a_5679_2511# a_3746_1779# a_5929_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1105 a_14494_13569# a_14407_13345# a_14090_13455# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1106 a_127_3207# a_9097_5098# a_10073_7110# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.325 pd=1.65 as=0.3 ps=2.6 w=1 l=0.15
X1107 a_3250_14835# a_2703_13747# a_3140_14835# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X1108 a_12174_11179# a_1225_10715# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1109 a_127_3207# a_3136_14540# a_3074_14657# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1110 w_62_10153# a_2371_10483# a_2539_10457# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1111 a_14323_2689# a_13541_2323# a_14239_2689# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1112 a_1229_14541# a_534_14471# a_1147_14541# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1113 w_62_361# a_13887_121# a_13835_147# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1114 a_127_3207# a_12231_8825# a_12179_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1115 w_62_10153# a_14368_11687# a_14407_11813# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1116 a_127_3207# a_13835_1235# a_15131_2145# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1117 a_2442_11571# a_2316_11687# a_2038_11703# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1118 a_11300_11571# a_11279_10695# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8 ad=0.9 pd=6.6 as=0.45 ps=3.3 w=3 l=0.15
X1119 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1120 a_127_3207# a_12854_9939# a_14125_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1121 a_727_15353# a_1147_14541# a_1397_14541# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1122 a_12231_7737# a_12402_7915# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X1123 a_13634_15599# a_14838_15701# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X1124 a_14708_513# a_14494_513# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1125 a_1147_13453# a_534_13383# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1126 a_14494_14657# a_14368_14559# a_14090_14543# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1127 a_127_3207# a_1783_147# a_3079_1057# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1128 a_905_2145# a_861_1753# a_739_2157# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1129 a_1208_1069# a_293_697# a_861_665# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1130 a_127_3207# a_3763_8825# a_5003_10189# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1131 a_2511_8000# a_2316_8031# a_2821_7763# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1132 a_15126_13569# a_14368_13471# a_14563_13440# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1133 a_14079_12300# div_out2_2 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1134 a_6185_3881# a_9585_3769# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X1135 a_14708_12659# a_14494_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1136 a_4137_7908# a_3660_7915# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1137 a_127_3207# a_2539_10207# a_2970_10261# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1138 a_1317_10803# a_1225_10715# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1139 a_127_3207# a_3746_9395# a_4575_10127# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1140 a_3136_1484# a_3250_1779# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X1141 a_12600_8673# a_12179_7763# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1142 a_3465_15407# a_1225_15531# a_3379_15407# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1143 a_1383_14051# a_1208_14125# a_1562_14113# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1144 a_127_3207# a_2371_15745# a_2539_15647# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1145 a_4711_11285# a_4077_12724# a_4137_12618# w_62_11241# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=1
X1146 a_12345_8313# a_12179_8313# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1147 a_861_11269# a_643_11027# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1148 a_127_3207# a_2371_10305# a_2539_10207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1149 a_1946_10483# a_1673_10489# a_1861_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1150 a_2511_9088# a_2355_8993# a_2656_9217# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1151 w_62_14505# a_1835_14265# a_1783_14291# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1152 a_2754_13979# a_941_13203# a_2880_14113# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1153 w_62_361# a_947_969# a_1835_121# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1154 a_12586_7943# a_13435_8611# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1155 a_12600_9761# a_12179_8851# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1156 a_2027_1753# div_fb3_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1157 a_127_3207# a_2316_11687# a_2355_11813# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1158 a_13541_9939# a_13375_9939# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1159 a_12600_15201# a_12179_14291# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1160 a_15126_11571# a_14407_11813# a_14563_11545# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1161 w_62_12329# a_12993_12659# a_14806_12267# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X1162 a_1225_10715# a_3660_12891# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1163 a_13814_10483# a_13541_10489# a_13729_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1164 a_127_3207# a_7331_4818# a_8109_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X1165 a_127_3207# a_122_11179# a_127_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1166 a_127_3207# a_1835_13177# a_1783_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1167 a_14708_11571# a_14494_11571# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1168 a_14368_1503# a_12174_923# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1169 a_13614_12115# a_12854_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1170 a_15289_10483# a_15123_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1171 a_535_15531# a_2027_13721# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1172 w_62_361# div_fb1_0 a_1229_397# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1173 a_127_3207# a_12271_10483# a_13375_10489# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1174 a_12854_15379# a_12271_15629# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1175 a_14465_14835# div_out3_3 w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1176 w_62_13417# a_14806_13979# a_15302_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X1177 w_62_14505# a_534_14471# a_476_14657# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X1178 a_127_3207# a_15188_11545# a_15126_11571# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1179 a_13199_8013# a_12586_7943# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1180 a_14494_12659# a_14407_12901# a_14090_12791# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1181 a_127_3207# a_2114_10051# a_2072_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1182 a_127_3207# a_12586_12899# a_12826_13025# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X1183 a_127_3207# a_15123_2323# a_15289_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1184 a_12957_9761# a_12913_9369# a_12791_9773# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1185 a_2316_12775# a_122_11179# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1186 a_127_3207# a_13435_12089# a_13369_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1187 a_12993_147# a_12402_299# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1188 a_4150_1032# a_4711_1571# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X1189 a_2038_399# a_2316_415# a_2272_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1190 w_62_12329# a_2754_12267# a_2703_12115# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1191 a_127_3207# a_446_399# a_397_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1192 w_62_2537# a_4575_2511# a_4533_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1193 a_1397_9101# div_fb0_1 w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1194 a_1673_15379# a_1507_15379# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1195 a_127_3207# a_4137_7908# a_4077_7948# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.3 ps=2.6 w=1 l=1
X1196 w_62_11241# div_fb3_2 a_2057_11277# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1197 a_5085_10189# a_2864_10189# a_5003_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1198 a_14109_8307# a_14079_8281# a_12403_10091# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X1199 w_62_9065# a_1208_9773# a_1383_9699# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1200 a_2038_11703# a_2355_11813# a_2313_11937# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1201 a_548_12115# a_127_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1202 a_12499_10715# a_13199_12659# a_13449_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1203 a_15302_13747# a_14806_13979# a_15131_14113# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1204 a_643_15213# a_293_14841# a_548_15201# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1205 a_127_3207# a_12174_923# a_12179_1785# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1206 a_127_3207# w_62_4713# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1207 a_127_3207# a_1783_8851# a_2027_9369# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1208 a_127_3207# a_2754_11179# a_2703_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1209 a_12695_8685# a_12179_8313# a_12600_8673# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1210 w_62_13417# a_861_13721# a_751_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1211 a_11296_9003# a_11658_8851# a_11300_9101# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1212 a_14090_14543# a_14407_14433# a_14365_14291# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1213 a_13435_15139# a_12854_15379# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1214 a_12600_2145# a_12179_1235# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1215 a_11382_11571# a_11296_11803# a_11300_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1216 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1217 a_15126_12659# a_14368_12775# a_14563_12633# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1218 a_14494_11571# a_14407_11813# a_14090_11703# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1219 a_12791_1069# a_12179_697# a_12695_1069# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1220 a_127_3207# a_3136_396# a_3074_513# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1221 a_397_1235# a_350_1387# a_179_1209# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1222 a_1383_2083# a_1208_2157# a_1562_2145# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1223 a_2072_9939# a_1673_9939# a_1946_10305# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1224 a_127_3207# a_12595_10457# a_12271_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1225 a_2371_2689# a_1507_2323# a_2114_2435# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1226 a_127_3207# a_5679_10127# a_5419_9913# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1227 w_62_2537# a_121_2297# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1228 a_12435_15629# a_12403_15531# a_12353_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X1229 a_5003_2573# a_2864_2573# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1230 a_11658_14291# a_11382_14291# a_11300_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1231 w_62_2537# a_1225_2475# a_11279_311# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X1232 a_127_3207# w_62_6889# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1233 a_3140_13747# a_1783_13203# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X1234 a_13449_1235# div_out0_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1235 a_5679_15567# a_3746_14835# a_5929_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1236 a_11279_311# a_5853_802# a_11279_649# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.225 pd=2.1 as=0.1125 ps=1.05 w=0.75 l=0.15
X1237 a_14563_1472# a_14407_1377# a_14708_1601# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1238 a_15131_1057# a_12993_147# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1239 a_4575_2511# a_4315_2297# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1240 a_12586_12899# a_13435_12089# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1241 a_127_3207# a_6422_11089# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X1242 a_127_3207# a_12854_15379# a_14125_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1243 a_1946_10483# a_1507_10489# a_1861_10483# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1244 a_12595_10457# a_13199_11571# a_13449_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1245 a_9097_5098# enb_0 w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1246 w_62_7977# a_14368_8031# a_14407_7905# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1247 a_12803_8307# a_12345_8313# a_12695_8685# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1248 a_2880_1057# a_1783_147# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X1249 a_2316_14559# a_122_13979# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1250 a_127_3207# w_62_4713# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1251 a_947_8585# a_403_10189# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1252 a_127_3207# a_2511_8000# a_2442_8129# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1253 w_62_13417# a_2754_13979# a_2703_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1254 w_62_13417# a_947_14025# a_2656_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1255 a_861_665# a_643_1069# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1256 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1257 a_751_9395# a_947_8585# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1258 a_1371_15353# a_11903_13203# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1259 a_15126_11571# a_14368_11687# a_14563_11545# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1260 a_1383_11001# a_947_11001# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1261 a_3746_691# a_3617_1387# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1262 a_13369_2157# a_12345_1785# a_13260_2157# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1263 a_14239_15745# a_13541_15379# a_13982_15491# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1264 w_62_361# a_12913_665# a_12803_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1265 w_62_1449# a_1208_2157# a_1383_2083# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1266 a_12913_1753# a_12695_2157# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1267 a_12854_9939# a_12271_10189# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1268 a_3657_10483# a_3379_10821# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1269 a_127_3207# w_62_5801# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1270 w_62_6889# a_127_3207# w_62_6889# w_62_6889# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1271 a_1946_2689# a_1507_2323# a_1861_2323# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1272 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1273 a_3250_9395# a_2703_8307# a_3140_9395# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X1274 a_127_3207# a_1783_14291# a_3079_15201# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1275 a_13814_10305# a_13375_9939# a_13729_9939# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1276 a_446_8015# a_350_9003# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1277 a_2749_13025# a_947_11001# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1278 a_3899_2573# a_3657_2323# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1279 a_3136_8012# a_3250_8307# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1280 a_14365_13025# a_13887_12633# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1281 a_12449_8851# a_12402_9003# a_12231_8825# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1282 a_11382_1235# a_11296_1387# a_11300_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1283 a_4315_15353# a_3899_15629# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1284 w_62_5801# a_127_3207# w_62_5801# w_62_5801# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1285 a_12586_14471# a_13435_15139# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1286 a_15289_9939# a_15123_9939# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1287 w_62_4713# a_127_3207# w_62_4713# w_62_4713# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1288 w_62_13417# a_947_14025# a_1835_13177# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1289 a_2442_8129# a_2316_8031# a_2038_8015# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1290 a_1673_15379# a_1507_15379# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1291 a_15289_2323# a_15123_2323# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1292 a_2313_147# a_1835_121# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1293 a_13634_10159# a_14838_10261# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1294 a_5085_10483# a_2864_10483# a_5003_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1295 a_127_3207# a_12231_1209# a_12179_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1296 w_62_10153# a_12271_10189# a_13375_9939# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1297 a_10437_4858# a_9567_4858# a_10073_5400# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.65 ps=2.65 w=2 l=0.5
X1298 a_14494_9217# a_14368_9119# a_14090_9103# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1299 w_62_6889# a_127_3207# w_62_6889# w_62_6889# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1300 a_12595_15353# a_12586_14471# a_13449_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X1301 a_12600_12115# a_12179_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1302 w_62_5801# a_127_3207# w_62_5801# w_62_5801# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1303 w_62_10153# a_3763_8825# a_5085_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1304 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1305 a_476_13569# a_446_13455# a_179_13177# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X1306 w_62_12329# a_1383_12089# a_1370_12481# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1307 a_12695_15213# a_12345_14841# a_12600_15201# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1308 a_14090_8015# a_14407_7905# a_14365_7763# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1309 a_13940_9939# a_13541_9939# a_13814_10305# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1310 a_12913_13721# a_12695_14125# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1311 w_62_10153# a_12586_9031# a_12528_9217# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X1312 w_62_10153# a_14755_8307# a_14806_9627# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X1313 a_127_3207# a_947_8585# a_905_9761# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1314 a_397_13025# a_534_12899# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1315 a_751_1779# a_947_969# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1316 a_5225_11511# a_4971_12724# a_4971_12724# w_62_11241# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1 as=0.15 ps=1.6 w=0.5 l=0.15
X1317 a_127_3207# a_3660_12891# a_5853_11873# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X1318 a_127_3207# a_14732_15629# a_15123_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1319 a_15126_9217# a_14368_9119# a_14563_9088# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1320 a_3140_8307# a_1783_7763# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X1321 a_12174_13979# a_1225_15531# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1322 a_15188_13452# a_15302_13747# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1323 a_13729_9939# a_13634_10159# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1324 a_774_7763# a_446_8015# a_350_7915# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1325 w_62_15593# a_2371_15745# a_2539_15647# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X1326 a_127_3207# a_13435_8611# a_13369_8685# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1327 a_2511_14528# a_2355_14433# a_2656_14657# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1328 a_14239_10305# a_13541_9939# a_13982_10051# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1329 a_127_3207# a_13199_12659# a_12499_10715# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1330 a_3250_1779# a_2703_691# a_3140_1779# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X1331 a_2073_13203# a_2038_13455# a_1835_13177# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1332 a_12600_1057# a_12179_147# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1333 a_15188_396# a_15302_691# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X1334 a_3074_8129# a_2316_8031# a_2511_8000# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1335 a_127_3207# a_6422_209# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=6
X1336 w_62_10153# a_12586_9031# a_13449_9101# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1337 a_12345_697# a_12179_697# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1338 a_9151_7110# a_9097_5098# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.105 pd=1.21 as=0.3 ps=2.6 w=1 l=0.15
X1339 a_3746_8307# a_3617_9003# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1340 w_62_15593# a_403_15629# a_1507_15379# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1341 a_5853_13858# a_3763_14265# a_5678_13470# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X1342 a_1861_2323# a_1766_2543# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1343 a_2821_8851# a_2442_9217# a_2749_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1344 a_14732_2573# a_14407_2591# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1345 a_127_3207# w_62_3625# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1346 w_62_12329# a_947_11001# a_2656_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1347 a_2114_10051# a_1946_10305# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1348 a_15131_14113# a_12993_13203# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1349 a_127_3207# a_6422_209# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X1350 a_11279_649# a_5853_802# a_11279_311# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.1125 pd=1.05 as=0.225 ps=2.1 w=0.75 l=0.15
X1351 a_2313_8851# a_1835_8825# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1352 w_62_2537# a_7331_5294# a_8109_6368# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X1353 a_1835_121# a_2038_399# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1354 a_14563_9088# a_14368_9119# a_14873_8851# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1355 w_62_14505# a_534_14471# a_1397_14541# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1356 a_4575_2511# a_3746_1779# a_4825_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1357 a_12296_4858# a_8169_4818# a_11749_5294# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.3 ps=2.6 w=1 l=0.15
X1358 a_13281_1485# a_12586_1415# a_13199_1485# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1359 a_293_1785# a_127_1785# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1360 a_127_3207# a_8169_4818# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=2
X1361 a_4077_12724# a_4077_12724# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X1362 a_127_3207# a_9097_5098# a_9887_7110# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.105 ps=1.21 w=1 l=0.15
X1363 a_127_3207# a_5419_15353# a_3763_14265# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1364 a_751_13747# a_947_14025# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1365 a_127_3207# a_11989_15353# a_12449_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1366 a_631_15531# a_534_13383# a_1397_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X1367 a_127_3207# a_13199_11571# a_12595_10457# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1368 w_62_2537# a_14755_691# a_14806_2011# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X1369 a_14109_691# a_13835_147# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1370 a_12957_2145# a_12913_1753# a_12791_2157# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1371 a_127_3207# a_2114_15491# a_2072_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1372 a_751_13747# a_293_13753# a_643_14125# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1373 a_6964_4858# a_6332_5146# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.32 as=0.33 ps=2.32 w=0.5 l=2.5
X1374 w_62_12329# a_947_11001# a_1835_12633# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1375 w_62_11241# a_947_11001# a_2656_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1376 a_13743_5587# a_6185_3209# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1377 a_127_3207# a_14239_10483# a_14407_10457# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1378 a_727_9913# a_534_9031# a_1397_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X1379 a_127_3207# a_1225_15531# a_5175_13488# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.075 ps=0.8 w=0.5 l=0.15
X1380 a_127_3207# a_6422_209# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X1381 a_127_3207# a_14732_2573# a_15123_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1382 a_122_923# a_1371_2297# a_1317_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1383 w_62_10153# a_14806_9627# a_15302_9395# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X1384 a_947_8585# a_403_10189# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1385 a_2272_513# a_1835_121# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1386 w_62_9065# a_2703_8307# a_2754_9627# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X1387 a_5637_10189# a_5003_10189# a_5419_9913# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1388 a_2057_14835# a_2027_14809# a_397_15531# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X1389 a_3899_15629# a_3657_15379# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1390 a_2371_15745# a_1507_15379# a_2114_15491# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1391 a_12803_13747# a_12854_15379# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1392 a_476_12659# a_446_12633# a_179_12633# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X1393 a_15302_14835# a_14755_13747# a_15192_14835# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X1394 a_127_3207# a_5679_10457# a_5419_10457# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1395 a_1229_9101# a_534_9031# a_1147_9101# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1396 a_2041_15745# a_1507_15379# a_1946_15745# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1397 a_739_14125# a_127_13753# a_643_14125# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1398 a_127_3207# a_1383_15139# a_1317_15213# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1399 w_62_10153# a_3763_11545# a_5085_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1400 w_62_12329# a_12913_12357# a_12803_12481# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1401 a_11296_11803# a_11658_11571# a_11300_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1402 w_62_10153# a_12174_11179# a_12179_11027# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1403 a_12528_13569# a_12498_13455# a_12231_13177# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X1404 a_127_3207# a_727_10457# a_403_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1405 a_127_3207# a_179_14265# a_127_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1406 a_13422_9395# a_12179_9401# a_13260_9773# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1407 a_12449_13025# a_12586_12899# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1408 w_62_2537# a_12586_1415# a_12402_1387# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X1409 a_127_3207# div_fb3_1 a_2245_9715# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1410 w_62_13417# div_out1_3 a_13281_13453# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1411 a_1208_15213# a_293_14841# a_861_14809# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1412 a_905_14113# a_861_13721# a_739_14125# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1413 a_1861_10483# a_1766_10647# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1414 w_62_10153# a_4575_10127# a_4533_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1415 a_127_3207# a_15123_10483# a_15289_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1416 w_62_11241# a_947_11001# a_1835_11545# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1417 w_62_13417# a_12586_13383# a_12528_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X1418 w_62_12329# div_fb1_2 a_1229_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1419 a_14806_9627# a_14755_8307# a_14932_9761# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1420 w_62_11241# a_3763_11545# a_3660_11179# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1421 a_3250_14835# a_2754_15067# a_3079_15201# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1422 a_127_3207# a_7331_4818# a_8109_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X1423 a_127_3207# a_2754_9627# a_2703_9395# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1424 a_13909_10305# a_13375_9939# a_13814_10305# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1425 a_12803_691# a_12345_697# a_12695_1069# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1426 w_62_15593# a_14407_15647# a_14323_15745# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1427 w_62_15593# a_2114_15491# a_2041_15745# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1428 a_1317_14125# a_293_13753# a_1208_14125# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1429 a_15188_1484# a_15302_1779# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1430 w_62_12329# a_2511_12633# a_2442_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1431 a_11279_649# enb_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X1432 a_14801_7763# a_12854_9939# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1433 a_127_3207# a_6422_13265# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=6
X1434 a_2754_8539# a_941_7763# a_2880_8673# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1435 a_127_3207# a_403_15629# a_1507_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1436 a_476_11571# a_121_10748# a_179_11545# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X1437 a_127_3207# a_1783_147# a_2027_665# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1438 a_15188_11545# a_15302_11393# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X1439 w_62_14505# a_1208_15213# a_1383_15139# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1440 a_12993_7763# a_12402_7915# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1441 a_3250_11393# a_2703_12115# a_3140_11393# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X1442 a_2038_399# a_2355_289# a_2313_147# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1443 a_13435_14051# a_13260_14125# a_13614_14113# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1444 a_631_2475# a_534_327# a_1397_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X1445 a_643_9773# a_293_9401# a_548_9761# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1446 a_13449_14291# div_out0_3 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1447 a_3074_8129# a_2355_7905# a_2511_8000# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1448 w_62_2537# a_14806_2011# a_15302_1779# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X1449 a_643_1069# a_127_697# a_548_1057# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1450 w_62_1449# a_2703_691# a_2754_2011# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X1451 a_5853_802# a_3746_691# a_5678_1571# w_62_1449# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X1452 a_12353_10189# a_12265_10091# a_12271_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X1453 a_14806_13979# a_12993_13203# a_14932_14113# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1454 a_3140_691# a_1783_147# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X1455 w_62_15593# a_13887_14265# a_13835_14291# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1456 w_62_361# a_3136_396# a_3074_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1457 a_3250_9395# a_2754_9627# a_3079_9761# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1458 a_2245_14067# a_1783_13203# a_535_15531# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X1459 a_127_3207# a_14368_11687# a_14407_11813# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1460 a_643_12115# a_293_12115# a_548_12115# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1461 w_62_11241# div_fb0_2 a_1229_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1462 a_13541_2323# a_13375_2323# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1463 a_947_969# a_403_2573# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1464 a_127_3207# w_62_4713# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1465 a_127_3207# a_1783_13203# a_2027_13721# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1466 a_13422_1779# a_12179_1785# a_13260_2157# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1467 a_8109_5400# a_6185_3881# a_8019_5400# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=0.15
X1468 a_127_3207# a_13887_7737# a_13835_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1469 w_62_11241# a_2511_11545# a_2442_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1470 a_11648_4958# enb_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X1471 a_127_3207# a_13887_13177# a_13835_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1472 a_2038_1487# a_2316_1503# a_2272_1601# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1473 a_127_3207# a_6422_13265# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X1474 a_12403_15531# a_14079_13721# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1475 a_12449_1235# a_12402_1387# a_12231_1209# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1476 w_62_2537# a_12183_5294# a_12183_5294# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=0.5
X1477 a_1229_397# a_534_327# a_1147_397# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1478 a_127_3207# a_3746_14835# a_4575_15567# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1479 a_5929_10189# a_5419_9913# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1480 w_62_361# a_4910_920# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X1481 a_12854_2323# a_12271_2573# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1482 a_127_3207# a_12854_9939# a_12957_8673# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1483 a_12803_13747# a_12345_13753# a_12695_14125# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1484 a_14079_9369# a_13835_8851# a_14465_9395# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1485 a_127_3207# a_13982_10051# a_13940_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1486 a_127_3207# a_4575_10127# a_4315_9913# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1487 a_947_11001# a_403_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1488 a_5637_10483# a_5003_10483# a_5419_10457# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1489 a_1317_9939# a_1225_10091# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1490 a_1397_14541# div_fb0_3 w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1491 a_6485_5594# a_6485_5594# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.33 pd=2.32 as=0.33 ps=2.32 w=0.5 l=3
X1492 a_2656_14657# a_2442_14657# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1493 a_14494_1601# a_14368_1503# a_14090_1487# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1494 w_62_10153# a_121_9913# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1495 a_14365_10861# a_13375_10489# a_14239_10483# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1496 a_2072_10861# a_1673_10489# a_1946_10483# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X1497 a_12528_12659# a_12498_12633# a_12231_12633# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X1498 a_397_147# a_350_299# a_179_121# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1499 a_11658_8851# a_11382_8851# a_11300_9101# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1500 a_15289_2323# a_15123_2323# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1501 a_127_3207# div_out3_0 a_14297_2099# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1502 a_12183_5294# a_10437_4858# a_12296_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.15 ps=1.3 w=1 l=0.15
X1503 a_127_3207# a_12174_11179# a_12179_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1504 w_62_4713# a_127_3207# w_62_4713# w_62_4713# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1505 a_548_8673# a_127_7763# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1506 a_127_3207# a_947_969# a_905_2145# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1507 a_12449_14291# a_12402_14443# a_12231_14265# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1508 a_1397_13203# div_fb1_3 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1509 a_127_3207# a_3660_13355# a_5853_13858# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X1510 a_2749_7763# a_947_8585# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1511 w_62_12329# a_12586_12899# a_12528_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X1512 a_13634_2543# a_14838_2645# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.154 ps=1.335 w=1 l=0.15
X1513 w_62_361# a_12854_2323# a_13887_121# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1514 a_127_3207# a_4315_10457# a_3617_11803# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1515 a_4711_1571# a_4077_332# a_4137_292# w_62_1449# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=1
X1516 w_62_10153# a_4575_10457# a_4533_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1517 a_1835_14265# a_2038_14543# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1518 a_127_3207# a_13435_995# a_13369_1069# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1519 a_12074_7210# a_7331_4818# a_7331_5294# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X1520 a_12265_10091# a_14079_9369# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1521 a_5085_15629# a_2864_15629# a_5003_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1522 a_127_3207# a_1835_121# a_1783_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1523 a_3657_2323# a_3379_2351# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1524 a_2027_8281# a_1783_7763# a_2413_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1525 w_62_5801# a_127_3207# w_62_5801# w_62_5801# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1526 a_127_3207# a_947_14025# a_905_14113# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1527 a_14239_2689# a_13375_2323# a_13982_2435# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1528 a_1208_14125# a_127_13753# a_861_13721# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1529 a_127_3207# a_3136_12633# a_3074_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1530 a_2754_12267# a_1783_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X1531 a_127_3207# a_14806_13979# a_14755_13747# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1532 a_1371_2297# a_11903_147# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1533 a_1766_2543# a_2970_2645# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1534 w_62_12329# a_941_12659# a_2754_12267# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X1535 a_127_3207# w_62_6889# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1536 w_62_10153# a_1371_9913# a_12174_8539# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1537 a_535_10091# a_2027_8281# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1538 a_2864_10189# a_2539_10207# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1539 a_1562_14113# a_947_14025# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1540 a_1766_10647# a_2970_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1541 a_127_3207# a_3136_9100# a_3074_9217# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1542 a_15192_13747# a_13835_13203# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X1543 a_2821_1235# a_2442_1601# a_2749_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1544 a_179_14265# a_350_14443# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X1545 a_12528_11571# a_11989_10748# a_12231_11545# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X1546 a_14079_1753# a_13835_1235# a_14465_1779# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1547 w_62_10153# div_out0_1 a_13281_9101# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1548 a_2313_1235# a_1835_1209# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1549 a_12345_14841# a_12179_14841# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1550 a_14563_1472# a_14368_1503# a_14873_1235# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1551 a_2442_14657# a_2355_14433# a_2038_14543# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1552 w_62_1449# a_3763_1209# a_3660_2011# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1553 w_62_7977# a_534_7943# a_350_7915# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X1554 w_62_9065# a_179_8825# a_127_8851# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X1555 a_12353_10483# a_12265_10715# a_12271_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X1556 w_62_10153# a_12586_11811# a_12528_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X1557 a_14090_399# a_14368_415# a_14324_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1558 a_14079_9369# div_out3_1 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1559 a_14708_9217# a_14494_9217# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1560 a_403_15629# a_631_15531# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X1561 a_15289_10483# a_15123_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1562 a_12695_12115# a_12345_12115# a_12600_12115# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1563 a_13435_11001# a_12854_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1564 a_13814_15745# a_13375_15379# a_13729_15379# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X1565 a_127_3207# div_out1_2 a_13199_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1566 a_1562_9761# a_947_8585# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1567 w_62_12329# a_2316_12775# a_2355_12901# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1568 a_127_3207# a_403_2573# a_1507_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1569 a_1229_12659# a_534_12899# a_1147_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1570 a_4273_2573# a_3899_2573# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1571 a_3660_11179# a_3617_11803# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1572 a_127_3207# a_12271_10189# a_13375_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1573 a_2656_8129# a_2442_8129# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1574 w_62_9065# a_5225_9261# a_5225_9261# w_62_9065# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.125 ps=1 w=0.5 l=0.15
X1575 a_2057_9395# a_1783_8851# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1576 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1577 a_12231_121# a_12402_299# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X1578 a_631_10715# a_1147_12659# a_1397_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1579 a_127_3207# a_13835_14291# a_15131_15201# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1580 a_5929_10483# a_5419_10457# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1581 a_2057_11277# a_1783_11571# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1582 w_62_361# a_1383_995# a_1370_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1583 a_13729_15379# a_13634_15599# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1584 a_631_2475# a_1147_397# a_1397_397# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1585 w_62_2537# a_14407_2591# a_14838_2645# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X1586 a_727_2297# a_534_1415# a_1397_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X1587 a_643_15213# a_127_14841# a_548_15201# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1588 a_3074_14657# a_2316_14559# a_2511_14528# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1589 w_62_15593# a_1225_15531# a_11279_13367# w_62_15593# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X1590 w_62_14505# a_5225_14701# a_5225_14701# w_62_14505# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.125 ps=1 w=0.5 l=0.15
X1591 a_2821_11937# a_2442_11571# a_2749_11937# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1592 a_14932_12115# a_13835_12659# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X1593 a_1383_8611# a_947_8585# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1594 a_1370_13747# a_127_13753# a_1208_14125# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1595 a_2027_11212# a_1783_11571# a_2413_11277# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1596 a_12791_15213# a_12179_14841# a_12695_15213# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1597 a_127_3207# a_727_9913# a_403_10189# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1598 a_127_3207# div_fb0_1 a_1147_9101# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1599 w_62_2537# a_14407_2591# a_14323_2689# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1600 w_62_13417# a_12854_15379# a_13887_13177# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1601 a_13982_2435# a_13814_2689# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1602 a_1835_8825# a_2038_9103# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1603 a_12271_10483# a_12499_10715# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X1604 a_127_3207# div_out0_2 a_13199_11571# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1605 a_1229_11571# a_534_11811# a_1147_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1606 w_62_1449# a_4077_332# a_5678_1571# w_62_1449# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X1607 w_62_10153# a_1225_10715# a_11279_10695# w_62_10153# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.15
X1608 a_727_10457# a_1147_11571# a_1397_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1609 a_534_327# a_1383_995# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1610 a_12345_1785# a_12179_1785# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1611 a_12695_8685# a_12345_8313# a_12600_8673# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1612 w_62_12329# a_1835_12633# a_1783_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1613 w_62_12329# a_13435_12089# a_13422_12481# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1614 a_12528_1601# a_11989_2297# a_12231_1209# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X1615 w_62_361# a_1208_1069# a_1383_995# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1616 a_14806_2011# a_14755_691# a_14932_2145# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1617 a_127_3207# a_6422_11089# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X1618 a_9193_6328# a_6332_6922# a_8019_6368# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.15 ps=1.3 w=1 l=0.5
X1619 a_179_8825# a_350_9003# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X1620 a_127_3207# div_out2_3 a_14297_14067# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1621 a_4711_14627# a_4077_13388# a_4137_13348# w_62_14505# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=1
X1622 a_8199_5400# a_8169_4818# a_8109_5400# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=0.15
X1623 a_127_3207# a_12854_15379# a_12957_14113# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1624 a_14563_13440# a_14368_13471# a_14873_13203# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1625 a_2497_9939# a_1507_9939# a_2371_10305# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X1626 a_127_3207# a_3617_14443# a_3899_15629# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1627 a_127_3207# a_2316_14559# a_2355_14433# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1628 a_127_3207# a_1147_9101# a_727_9913# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1629 w_62_15593# a_3763_14265# a_5085_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1630 w_62_14505# a_2754_15067# a_3250_14835# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X1631 a_2057_1779# a_1783_1235# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1632 a_2316_13471# a_122_13979# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1633 a_2754_923# a_941_147# a_2880_1057# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1634 w_62_1449# a_5225_1645# a_5225_1645# w_62_1449# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.125 ps=1 w=0.5 l=0.15
X1635 a_127_3207# a_11648_4958# a_11648_4958# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=0.5
X1636 w_62_10153# a_1371_10457# a_12174_11179# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1637 a_14563_14528# a_14407_14433# a_14708_14657# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X1638 a_127_3207# a_446_13455# a_397_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1639 a_14806_15067# a_13835_14291# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X1640 a_2864_10483# a_2539_10457# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1641 a_14324_9217# a_13887_8825# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1642 a_14125_13203# a_14090_13455# a_13887_13177# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1643 a_14368_11687# a_12174_11179# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1644 a_643_2157# a_293_1785# a_548_2145# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1645 a_127_3207# a_15188_14540# a_15126_14657# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1646 a_13281_14541# a_12586_14471# a_13199_14541# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1647 a_127_3207# div_fb2_0 a_2245_1011# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1648 a_2272_8129# a_1835_7737# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1649 w_62_15593# a_12854_15379# a_14708_14657# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1650 w_62_10153# a_14806_11179# a_14755_11027# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1651 a_350_1387# a_121_2297# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X1652 a_14125_7763# a_14090_8015# a_13887_7737# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X1653 a_12127_10133# a_127_3207# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1654 a_5419_9913# a_5003_10189# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1655 a_127_3207# a_2539_10207# a_2497_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1656 w_62_2537# a_13887_1209# a_13835_1235# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1657 a_127_3207# a_2511_12633# a_2442_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1658 a_14494_11571# a_14368_11687# a_14090_11703# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1659 a_12600_11027# a_12179_11571# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1660 a_12402_7915# a_12498_8015# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X1661 a_293_9401# a_127_9401# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1662 w_62_11241# a_1835_11545# a_1783_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1663 a_3250_1779# a_2754_2011# a_3079_2145# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1664 a_127_3207# a_1147_13453# a_631_15531# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1665 a_739_11027# a_127_11027# a_643_11027# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1666 a_4971_13388# a_4137_13348# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X1667 a_127_3207# a_13835_12659# a_14079_12300# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1668 a_127_3207# a_2754_923# a_2703_691# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1669 a_2316_8031# a_122_8539# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1670 a_2316_9119# a_122_8539# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1671 a_13199_13453# a_12586_13383# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1672 a_3617_14443# a_3899_15629# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1673 a_11279_8265# a_3660_7915# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X1674 w_62_2537# a_12271_2573# a_13375_2323# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1675 a_13449_8013# div_out1_1 w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1676 w_62_7977# a_1383_8611# a_1370_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1677 a_127_3207# a_3519_15381# a_3465_15407# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1678 a_2864_15629# a_2539_15647# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1679 a_127_3207# a_12854_2323# a_12957_1057# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X1680 a_2316_12775# a_122_11179# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1681 a_127_3207# a_3660_13355# a_11296_14443# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X1682 a_122_13979# a_1371_15353# a_1317_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1683 a_127_3207# a_4137_12618# a_4077_12724# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.3 ps=2.6 w=1 l=1
X1684 w_62_11241# a_1225_10715# a_4971_12724# w_62_11241# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1 as=0.15 ps=1.6 w=0.5 l=0.15
X1685 w_62_2537# a_7331_5294# a_7331_4818# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X1686 a_12695_15213# a_12179_14841# a_12600_15201# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1687 a_127_3207# a_13835_7763# a_14079_8281# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1688 w_62_12329# a_12854_10483# a_13887_12633# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1689 a_10073_5400# enb_0 w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.65 ps=2.65 w=2 l=0.15
X1690 a_127_3207# a_1783_8851# a_3079_9761# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1691 a_127_3207# a_3519_9941# a_3465_9967# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X1692 a_1317_11027# a_293_11027# a_1208_11027# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1693 a_12913_11269# a_12695_11027# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1694 a_2442_1601# a_2355_1377# a_2038_1487# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1695 a_643_9773# a_127_9401# a_548_9761# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1696 a_293_12115# a_127_12115# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1697 a_1371_15353# a_11903_13203# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1698 a_12174_923# a_1371_2297# a_13185_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1699 a_6485_6328# a_6485_6328# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.33 pd=2.32 as=0.33 ps=2.32 w=0.5 l=3
X1700 a_403_2573# a_631_2475# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X1701 a_1861_2323# a_1766_2543# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X1702 a_14109_14835# a_14079_14809# a_12265_15531# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X1703 a_6185_3321# a_9567_6368# a_10073_6368# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.65 ps=2.65 w=2 l=0.5
X1704 a_2027_14809# div_fb3_3 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1705 a_1371_10457# a_11903_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X1706 a_3074_513# a_2355_289# a_2511_384# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1707 w_62_10153# a_14806_9627# a_14755_9395# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1708 w_62_2537# a_12854_2323# a_14708_1601# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1709 a_127_3207# a_12586_327# a_12826_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X1710 w_62_3625# a_127_3207# w_62_3625# w_62_3625# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1711 a_14079_14809# a_13835_14291# a_14465_14835# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1712 a_127_3207# w_62_4713# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1713 w_62_7977# a_13260_8685# a_13435_8611# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1714 a_122_923# a_1225_2475# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1715 a_127_3207# a_534_7943# a_774_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X1716 a_12803_8307# a_12854_9939# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X1717 a_12271_2573# a_12499_2475# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X1718 a_947_14025# a_403_15629# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1719 a_127_3207# a_15123_15379# a_15289_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1720 a_5637_15629# a_5003_15629# a_5419_15353# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1721 w_62_10153# a_12854_9939# a_13887_8825# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1722 w_62_9065# a_1835_8825# a_1783_8851# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1723 w_62_11241# a_4077_12724# a_5678_11285# w_62_11241# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X1724 w_62_4713# a_127_3207# w_62_4713# w_62_4713# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1725 a_1397_7763# div_fb1_1 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1726 a_751_9395# a_293_9401# a_643_9773# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1727 w_62_10153# a_12854_10483# a_13887_11545# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1728 w_62_361# a_12586_327# a_13449_397# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1729 a_534_9031# a_1383_9699# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1730 w_62_7977# a_947_8585# a_1835_7737# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1731 w_62_7977# div_fb2_1 a_2057_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1732 a_127_3207# a_3136_1484# a_3074_1601# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X1733 a_5853_11873# a_6422_11089# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X1734 w_62_1449# a_3136_1484# a_3074_1601# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1735 a_548_15201# a_127_14291# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1736 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1737 a_127_3207# a_4315_9913# a_3617_9003# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1738 a_1371_2297# a_11903_147# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X1739 w_62_7977# a_12231_7737# a_12179_7763# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X1740 w_62_12329# a_14563_12633# a_14494_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1741 w_62_10153# div_out3_2 a_14109_11277# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1742 w_62_15593# a_4575_15567# a_4533_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1743 w_62_7977# a_2754_8539# a_2703_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1744 a_446_13455# a_350_14443# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1745 a_14090_11703# a_14407_11813# a_14365_11937# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1746 w_62_4713# a_127_3207# w_62_4713# w_62_4713# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X1747 w_62_15593# a_13260_15213# a_13435_15139# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1748 a_127_3207# a_12231_14265# a_12179_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1749 a_643_2157# a_127_1785# a_548_2145# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1750 a_15302_11393# a_14755_12115# a_15192_11393# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X1751 a_12449_8851# a_12586_9031# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1752 w_62_9065# a_122_8539# a_127_9401# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1753 a_1397_147# div_fb1_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1754 a_14324_513# a_13887_121# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1755 a_476_8129# a_446_8015# a_179_7737# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X1756 w_62_361# a_2316_415# a_2355_289# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1757 w_62_2537# a_11279_311# a_11279_311# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.3 as=0.9 ps=6.6 w=3 l=0.15
X1758 a_12403_2475# a_14079_665# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1759 a_1317_8685# a_293_8313# a_1208_8685# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1760 w_62_15593# a_13982_15491# a_13909_15745# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1761 a_12957_12115# a_12913_12357# a_12791_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X1762 a_1562_2145# a_947_969# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1763 a_14801_13203# a_12854_15379# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X1764 a_14297_9715# a_13835_8851# a_12265_10091# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X1765 w_62_2537# a_14806_2011# a_14755_1779# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X1766 a_1208_11027# a_293_11027# a_861_11269# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1767 a_127_3207# a_1783_11571# a_3079_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1768 a_14297_14067# a_13835_13203# a_12403_15531# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X1769 a_14090_8015# a_14368_8031# a_14324_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X1770 a_3136_12633# a_3250_12481# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1771 a_127_3207# a_8169_4818# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=2
X1772 w_62_9065# a_2511_9088# a_2442_9217# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1773 a_13982_10457# a_13814_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X1774 w_62_361# a_12231_121# a_12179_147# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X1775 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1776 a_12913_8281# a_12695_8685# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1777 a_12345_697# a_12179_697# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1778 a_127_3207# a_5419_2297# a_3763_1209# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1779 a_13260_8685# a_12179_8313# a_12913_8281# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1780 a_14563_12633# a_14368_12775# a_14873_13025# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1781 a_127_3207# w_62_6889# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X1782 a_2245_8627# a_1783_7763# a_535_10091# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X1783 a_12353_15629# a_12265_15531# a_12271_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.13 pd=1.26 as=0.26 ps=2.52 w=1 l=0.15
X1784 a_2114_10457# a_1946_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X1785 a_397_13203# a_350_13355# a_179_13177# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1786 a_15302_8307# a_12993_7763# a_15192_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X1787 a_10437_4858# a_9567_4858# a_10073_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.325 ps=1.65 w=1 l=0.5
X1788 w_62_10153# a_14563_11545# a_14494_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1789 a_1370_691# a_127_697# a_1208_1069# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1790 a_1208_11027# a_127_11027# a_861_11269# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1791 w_62_1449# a_947_969# a_2656_1601# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X1792 a_751_1779# a_293_1785# a_643_2157# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X1793 a_534_1415# a_1383_2083# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1794 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1795 a_12791_9773# a_12179_9401# a_12695_9773# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1796 a_14079_665# div_out2_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1797 a_127_3207# a_13982_10457# a_13940_10861# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X1798 a_293_12115# a_127_12115# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1799 a_12231_13177# a_12402_13355# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X1800 a_127_3207# div_fb0_0 a_1147_1485# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1801 a_3465_2351# a_1225_2475# a_3379_2351# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1802 w_62_2537# enb_0 a_10073_5400# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.65 pd=2.65 as=0.6 ps=4.6 w=2 l=0.15
X1803 w_62_11241# a_1208_11027# a_1383_11001# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1804 a_403_10483# a_397_10715# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
X1805 a_127_3207# a_11279_12307# a_11279_12307# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.225 pd=1.8 as=0.45 ps=3.6 w=1.5 l=0.15
X1806 a_2754_923# a_1783_147# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X1807 a_127_3207# a_12498_12633# a_12449_13025# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1808 w_62_2537# a_3617_1387# a_3981_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1809 a_1225_15531# a_3660_13355# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1810 a_4137_13348# a_3660_13355# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X1811 a_14806_9627# a_13835_8851# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X1812 a_5929_15629# a_5419_15353# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1813 a_14708_14657# a_14494_14657# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X1814 a_13260_8685# a_12345_8313# a_12913_8281# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1815 a_3079_15201# a_2703_13747# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1816 a_15131_9761# a_14755_8307# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1817 a_127_3207# a_6422_7825# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X1818 a_941_7763# a_350_7915# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1819 a_2880_15201# a_1783_14291# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X1820 w_62_13417# a_12586_13383# a_13449_13453# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1821 a_12695_1069# a_12345_697# a_12600_1057# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X1822 w_62_2537# a_727_2297# a_673_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1823 a_3136_14540# a_3250_14835# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X1824 a_2880_9761# a_1783_8851# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X1825 w_62_12329# a_534_12899# a_1397_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1826 a_1383_995# a_947_969# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X1827 a_15192_691# a_13835_147# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X1828 a_3079_8673# a_941_7763# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1829 a_14873_7763# a_14494_8129# a_14801_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1830 a_1317_15379# a_1225_15531# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1831 w_62_361# a_15188_396# a_15126_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X1832 a_2413_12365# div_fb2_2 w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1833 a_127_3207# a_1147_1485# a_727_2297# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1834 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1835 w_62_7977# a_861_8281# a_751_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1836 a_127_3207# a_535_10715# a_403_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X1837 a_14365_7763# a_13887_7737# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1838 w_62_1449# a_2511_1472# a_2442_1601# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X1839 a_774_13203# a_446_13455# a_350_13355# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1840 w_62_12329# a_122_11179# a_127_12115# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1841 a_941_147# a_350_299# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1842 a_12499_2475# a_13199_397# a_13449_397# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X1843 a_2027_11212# div_fb3_2 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1844 a_3617_1387# a_3899_2573# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1845 a_2754_8539# a_1783_7763# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X1846 a_13614_14113# a_12854_15379# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X1847 a_127_3207# div_fb3_3 a_2245_15155# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1848 a_12498_13455# a_12402_14443# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1849 a_2442_513# a_2355_289# a_2038_399# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1850 a_4077_13388# a_4077_13388# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X1851 a_293_1785# a_127_1785# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1852 a_12791_12115# a_12179_12115# a_12695_12115# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1853 a_127_3207# a_2316_415# a_2355_289# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1854 a_14494_14657# a_14407_14433# a_14090_14543# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1855 w_62_11241# a_534_11811# a_1397_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1856 a_15289_15379# a_15123_15379# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1857 a_127_3207# a_446_8015# a_397_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X1858 w_62_15593# a_1371_15353# a_12174_13979# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1859 a_2313_11937# a_1835_11545# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X1860 a_13634_10647# a_14838_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X1861 a_2864_15629# a_2539_15647# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1862 a_2442_13569# a_2316_13471# a_2038_13455# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X1863 a_127_3207# a_6422_13265# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=6
X1864 a_127_3207# a_13435_14051# a_13369_14125# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1865 a_14806_2011# a_13835_1235# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X1866 a_127_3207# a_14563_384# a_14494_513# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X1867 a_5637_2573# a_5003_2573# a_5419_2297# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X1868 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1869 a_12499_10091# a_12586_7943# a_13449_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X1870 a_3746_1779# a_3660_2011# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1871 a_127_3207# a_5853_13858# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=3.3 pd=22.6 as=0 ps=0 w=11 l=2
X1872 a_14239_10483# a_13541_10489# a_13982_10457# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X1873 a_14873_13203# a_14494_13569# a_14801_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X1874 a_127_3207# a_3746_1779# a_5679_2511# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1875 w_62_12329# a_14368_12775# a_14407_12901# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1876 a_14465_8307# div_out2_1 w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1877 a_13260_14125# a_12345_13753# a_12913_13721# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1878 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X1879 a_8109_6368# a_6185_3321# a_8019_6368# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=0.15
X1880 a_12600_1057# a_12179_147# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X1881 a_1861_10483# a_1766_10647# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X1882 a_127_3207# a_12854_9939# a_14125_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1883 a_127_3207# a_947_11001# a_2073_11937# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1884 a_12231_8825# a_12402_9003# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X1885 a_11749_5294# a_12183_5294# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=0.5
X1886 a_12231_12633# a_12402_12891# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X1887 a_12913_11269# a_12695_11027# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1888 a_127_3207# a_1783_1235# a_3079_2145# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1889 a_2413_13747# div_fb2_3 w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1890 a_4137_13348# a_4137_13348# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.15 ps=1.3 w=1 l=1
X1891 a_14109_11277# a_13835_11571# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1892 a_127_3207# a_13887_121# a_13835_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X1893 a_127_3207# a_947_8585# a_2073_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X1894 a_15126_14657# a_14368_14559# a_14563_14528# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X1895 a_2511_9088# a_2316_9119# a_2821_8851# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X1896 a_259_15573# a_127_3207# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X1897 a_127_3207# a_1383_11001# a_1317_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X1898 a_13422_13747# a_12179_13753# a_13260_14125# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X1899 a_127_3207# a_14407_10207# a_14838_10261# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1900 a_127_3207# a_6422_13265# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X1901 w_62_10153# a_2539_10207# a_2970_10261# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X1902 a_1946_2689# a_1673_2323# a_1861_2323# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X1903 a_1397_1485# div_fb0_0 w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1904 a_12600_9761# a_12179_8851# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X1905 a_1383_15139# a_1208_15213# a_1562_15201# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X1906 a_11300_1485# a_11279_311# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.9 pd=6.6 as=0.45 ps=3.3 w=3 l=0.15
X1907 a_127_3207# a_12595_15353# a_12271_15629# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1908 a_127_3207# a_14407_15647# a_14365_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X1909 a_127_3207# a_14806_8539# a_14755_8307# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1910 a_12345_9401# a_12179_9401# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1911 a_861_12357# a_643_12115# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X1912 a_15126_13569# a_14407_13345# a_14563_13440# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X1913 a_9887_7110# a_9193_6328# a_8199_6368# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.105 pd=1.21 as=0.15 ps=1.3 w=1 l=0.5
X1914 a_4077_332# a_1225_2475# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.125 ps=1 w=0.5 l=0.15
X1915 w_62_13417# a_179_13177# a_127_13203# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X1916 a_2754_15067# a_2703_13747# a_2880_15201# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X1917 a_14368_415# a_12174_923# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1918 a_12586_9031# a_13435_9699# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1919 a_11658_11571# a_11382_11571# a_11300_11891# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X1920 a_12231_11545# a_12402_11803# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X1921 w_62_1449# a_534_1415# a_476_1601# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X1922 a_11296_1387# a_11658_1235# a_11300_1485# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X1923 a_3250_11393# a_2754_11179# a_3079_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1924 w_62_12329# a_13887_12633# a_13835_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1925 a_14732_10483# a_14407_10457# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1926 a_3465_10821# a_1225_10715# a_3379_10821# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X1927 a_2371_10483# a_1507_10489# a_2114_10457# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X1928 a_534_7943# a_1383_8611# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1929 a_127_3207# a_122_11179# a_127_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1930 a_127_3207# a_11279_13705# a_11279_13705# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.225 pd=1.8 as=0.45 ps=3.6 w=1.5 l=0.15
X1931 a_12826_13203# a_12498_13455# a_12402_13355# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X1932 a_1147_8013# a_534_7943# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1933 a_2455_15745# a_1673_15379# a_2371_15745# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1934 a_643_11027# a_127_11027# a_548_11027# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X1935 a_127_3207# a_14368_14559# a_14407_14433# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1936 a_5853_11873# a_3763_11545# a_5678_12642# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X1937 a_12074_7210# a_7331_4818# a_7331_5294# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X1938 a_397_15531# a_2027_14809# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X1939 w_62_15593# a_14806_15067# a_15302_14835# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X1940 a_2041_10483# a_1507_10489# a_1946_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X1941 a_12449_13025# a_12402_12891# a_12231_12633# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X1942 a_127_3207# a_534_13383# a_774_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X1943 w_62_7977# a_12174_8539# a_12179_8313# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1944 a_13199_9101# a_12586_9031# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1945 a_861_9369# a_643_9773# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X1946 a_12345_11027# a_12179_11027# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1947 a_14732_2573# a_14407_2591# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X1948 w_62_361# a_13435_995# a_13422_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X1949 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1950 a_3660_9627# a_3617_9003# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X1951 a_12449_1235# a_12586_1415# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1952 a_1317_1069# a_293_697# a_1208_1069# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X1953 a_14323_15745# a_13541_15379# a_14239_15745# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X1954 a_13449_13453# div_out1_3 w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1955 a_127_3207# a_2539_10457# a_2970_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X1956 a_8109_4858# a_6185_3881# a_8019_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.3 ps=2.6 w=1 l=0.15
X1957 a_127_3207# div_fb1_0 a_1147_397# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1958 a_3617_1387# a_4315_2297# a_4273_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X1959 a_3657_15379# a_3379_15407# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.182 pd=1.86 as=0.1118 ps=1.04 w=0.65 l=0.15
X1960 a_2038_13455# a_2355_13345# a_2313_13203# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X1961 a_127_3207# w_62_4713# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1962 a_127_3207# enb_0 a_5853_802# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X1963 a_12499_10715# a_12586_12899# a_13449_12979# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X1964 a_15192_9395# a_13835_8851# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X1965 a_1397_12659# div_fb1_2 w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1966 w_62_10153# a_13887_11545# a_13835_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X1967 w_62_12329# div_fb2_2 a_2057_12365# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X1968 a_127_3207# a_13199_13453# a_12499_15531# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.208 pd=1.94 as=0.25025 ps=1.42 w=0.65 l=0.15
X1969 w_62_10153# a_14407_10457# a_14323_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X1970 a_534_13383# a_1383_14051# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X1971 w_62_10153# a_2114_10457# a_2041_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X1972 a_13260_1069# a_12179_697# a_12913_665# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X1973 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X1974 a_15302_14835# a_14806_15067# a_15131_15201# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X1975 w_62_361# a_12174_923# a_12179_697# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X1976 a_293_13753# a_127_13753# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1977 a_127_3207# w_62_5801# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1978 a_5679_10127# a_5419_9913# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X1979 a_127_3207# a_2754_12267# a_2703_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X1980 a_1208_9773# a_293_9401# a_861_9369# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X1981 w_62_14505# a_861_14809# a_751_14835# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1982 a_13887_13177# a_14090_13455# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X1983 a_127_3207# a_3746_11027# a_5679_10457# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X1984 a_12586_327# a_13435_995# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X1985 a_127_3207# w_62_6889# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1986 w_62_11241# a_2754_11179# a_3250_11393# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X1987 a_2057_8307# a_2027_8281# a_535_10091# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X1988 w_62_13417# a_12993_13203# a_14806_13979# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X1989 a_14494_8129# a_14407_7905# a_14090_8015# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X1990 a_127_3207# div_fb3_2 a_2245_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X1991 w_62_361# a_13260_1069# a_13435_995# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X1992 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1993 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X1994 a_12791_2157# a_12179_1785# a_12695_2157# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X1995 a_14806_11179# a_13835_11571# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X1996 a_446_399# a_350_1387# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X1997 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X1998 w_62_361# a_861_665# a_751_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X1999 a_127_3207# a_122_8539# a_127_8313# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2000 a_11279_12307# a_3660_12891# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X2001 a_6185_3321# a_9585_3321# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X2002 a_12595_10457# a_12586_11811# a_13449_11891# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2003 a_14297_1011# a_13835_147# a_12403_2475# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X2004 a_3140_14835# a_1783_14291# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X2005 a_14368_11687# a_12174_11179# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2006 a_1397_11571# div_fb0_2 w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2007 a_861_1753# a_643_2157# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2008 a_15131_2145# a_14755_691# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2009 a_2272_13569# a_1835_13177# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2010 a_10437_4858# a_6185_3881# sky130_fd_pr__cap_mim_m3_1 l=7 w=7
X2011 a_2442_12659# a_2316_12775# a_2038_12791# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2012 w_62_10153# a_14368_9119# a_14407_8993# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2013 a_127_3207# a_14368_8031# a_14407_7905# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2014 w_62_13417# a_2316_13471# a_2355_13345# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2015 a_2511_1472# a_2355_1377# a_2656_1601# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2016 a_2880_2145# a_1783_1235# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X2017 a_3079_1057# a_941_147# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2018 a_14368_415# a_12174_923# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2019 a_8199_6368# a_6332_6922# a_9567_6368# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.3 ps=2.6 w=1 l=0.5
X2020 a_127_3207# w_62_5801# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2021 a_15192_1779# a_13835_1235# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X2022 w_62_6889# a_127_3207# w_62_6889# w_62_6889# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2023 a_127_3207# a_2511_9088# a_2442_9217# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2024 w_62_14505# a_947_14025# a_2656_14657# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1092 ps=1.36 w=0.42 l=0.15
X2025 w_62_14505# a_2754_15067# a_2703_14835# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2026 a_861_1753# a_643_2157# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2027 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2028 w_62_7977# a_2316_8031# a_2355_7905# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2029 a_548_14113# a_127_13203# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2030 a_1383_12089# a_947_11001# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2031 a_8199_6368# a_5853_802# a_8109_6368# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=0.15
X2032 w_62_7977# a_15188_8012# a_15126_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2033 a_350_299# a_446_399# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X2034 a_2371_2689# a_1673_2323# a_2114_2435# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2035 w_62_7977# a_534_7943# a_1397_8013# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2036 w_62_13417# div_fb2_3 a_2057_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2037 a_127_3207# a_6422_7825# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X2038 a_127_3207# a_4137_13348# a_5678_13470# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X2039 a_13449_397# div_out1_0 w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2040 a_12695_11027# a_12179_11027# a_12600_11027# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2041 a_14239_10305# a_13375_9939# a_13982_10051# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1095 ps=1.075 w=0.42 l=0.15
X2042 a_1208_2157# a_293_1785# a_861_1753# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2043 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2044 a_9151_5400# enb_0 w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.21 pd=2.21 as=0.6 ps=4.6 w=2 l=0.15
X2045 a_127_3207# a_12586_13383# a_12826_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X2046 a_12345_11027# a_12179_11027# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2047 a_2413_9395# div_fb3_1 w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2048 a_5853_8418# a_6422_7825# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X2049 a_2864_10189# a_2539_10207# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2050 a_1225_10091# a_3660_7915# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2051 w_62_2537# a_12586_1415# a_13449_1485# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2052 a_3136_9100# a_3250_9395# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2053 w_62_6889# a_127_3207# w_62_6889# w_62_6889# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2054 a_127_3207# a_1783_1235# a_2027_1753# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2055 a_1371_10457# a_11903_12659# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2056 w_62_5801# a_127_3207# w_62_5801# w_62_5801# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2057 w_62_14505# a_947_14025# a_1835_14265# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2058 a_127_3207# a_2316_12775# a_2355_12901# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2059 a_2442_9217# a_2316_9119# a_2038_9103# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2060 a_15126_12659# a_14407_12901# a_14563_12633# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2061 w_62_2537# enb_0 a_9887_5400# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.21 ps=2.21 w=2 l=0.15
X2062 a_2821_14291# a_2442_14657# a_2749_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2063 a_3746_13747# a_3617_14443# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2064 a_127_3207# a_179_12633# a_127_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2065 a_2038_8015# a_2355_7905# a_2313_7763# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2066 a_14873_147# a_14494_513# a_14801_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2067 a_13185_10803# a_1225_10715# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2068 a_13887_12633# a_14090_12791# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2069 a_127_3207# a_12854_2323# a_14125_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2070 a_6964_6922# a_6332_6922# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.33 pd=2.32 as=0.33 ps=2.32 w=0.5 l=2.5
X2071 a_397_10715# a_2027_11212# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X2072 a_127_3207# a_14239_15745# a_14407_15647# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2073 a_13260_14125# a_12179_13753# a_12913_13721# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2074 a_127_3207# a_13835_11571# a_15131_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2075 a_127_3207# a_15188_12633# a_15126_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2076 a_127_3207# div_out1_1 a_13199_8013# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2077 a_476_14657# a_121_15353# a_179_14265# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X2078 a_861_12357# a_643_12115# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2079 a_14090_9103# a_14407_8993# a_14365_8851# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2080 a_12913_14809# a_12695_15213# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2081 a_861_13721# a_643_14125# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2082 a_13887_7737# a_14090_8015# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2083 a_15289_2323# a_15123_2323# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2084 a_14109_8307# a_13835_7763# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2085 w_62_7977# a_12913_8281# a_12803_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2086 a_127_3207# a_4137_12618# a_5678_12642# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X2087 a_127_3207# a_179_7737# a_127_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2088 a_1371_9913# a_11903_7763# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2089 a_534_11811# a_1383_11001# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2090 a_15188_14540# a_15302_14835# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2091 a_2511_1472# a_2316_1503# a_2821_1235# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2092 a_127_3207# a_5679_15567# a_5419_15353# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2093 a_10073_6368# enb_0 w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.65 ps=2.65 w=2 l=0.15
X2094 a_739_8685# a_127_8313# a_643_8685# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2095 a_774_8851# a_121_9913# a_350_9003# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2096 a_127_3207# a_3617_9003# a_3899_10189# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2097 a_127_3207# a_13435_9699# a_13369_9773# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2098 a_127_3207# w_62_3625# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2099 a_2272_12659# a_1835_12633# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2100 a_11630_6516# a_7331_4818# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2101 a_127_3207# a_727_15353# a_403_15629# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2102 w_62_10153# a_13260_11027# a_13435_11001# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2103 a_12600_2145# a_12179_1235# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2104 a_3074_9217# a_2316_9119# a_2511_9088# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2105 a_13449_12979# div_out1_2 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2106 a_1225_2475# enb_0 w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2107 a_2413_1779# div_fb3_0 w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2108 a_2038_12791# a_2355_12901# a_2313_13025# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2109 a_127_3207# a_179_11545# a_127_11571# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2110 a_12345_1785# a_12179_1785# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2111 a_8199_4858# a_8169_4818# a_8109_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.15 ps=1.3 w=1 l=0.15
X2112 a_3074_14657# a_2355_14433# a_2511_14528# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2113 a_476_513# a_446_399# a_179_121# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X2114 a_127_3207# a_15123_15379# a_15289_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2115 a_13887_11545# a_14090_11703# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2116 w_62_9065# a_1225_10091# a_4971_7948# w_62_9065# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1 as=0.15 ps=1.6 w=0.5 l=0.15
X2117 a_127_3207# a_14563_11545# a_14494_11571# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2118 a_1229_1485# a_534_1415# a_1147_1485# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2119 a_13281_12659# a_12586_12899# a_13199_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2120 a_127_3207# a_12498_8015# a_12449_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2121 a_4137_12618# a_4077_12724# a_4711_11285# w_62_11241# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=1
X2122 a_15131_15201# a_14755_13747# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2123 a_13729_10483# a_13634_10647# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2124 w_62_13417# a_122_13979# a_127_13753# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2125 a_12854_9939# a_12271_10189# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2126 w_62_361# a_14368_415# a_14407_289# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2127 a_127_3207# enb_0 a_11296_1387# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X2128 a_5679_10457# a_5419_10457# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2129 a_2455_2689# a_1673_2323# a_2371_2689# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2130 a_2511_14528# a_2316_14559# a_2821_14291# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2131 a_127_3207# a_3763_1209# a_5003_2573# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2132 a_12600_14113# a_12179_13203# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2133 a_12499_10091# a_13199_8013# a_13449_8013# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X2134 w_62_13417# a_1383_14051# a_1370_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2135 a_13940_15379# a_13541_15379# a_13814_15745# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2136 a_11279_13705# a_5853_13858# a_11279_13367# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.1125 pd=1.05 as=0.225 ps=2.1 w=0.75 l=0.15
X2137 a_13541_15379# a_13375_15379# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2138 a_751_14835# a_947_14025# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2139 a_127_3207# a_2539_2591# a_2970_2645# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2140 a_2749_13203# a_947_14025# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2141 a_2272_11571# a_1835_11545# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2142 a_127_3207# a_3746_1779# a_4575_2511# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2143 a_14365_13203# a_13887_13177# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2144 a_13449_11891# div_out0_2 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2145 a_13199_1485# a_12586_1415# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2146 a_3660_9627# a_3763_8825# a_3709_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2147 a_14368_8031# a_12174_8539# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2148 a_13422_691# a_12179_697# a_13260_1069# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2149 a_127_3207# a_2371_2689# a_2539_2591# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2150 w_62_10153# a_3617_9003# a_3981_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2151 a_11382_14291# a_11296_14443# a_11300_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2152 a_751_14835# a_293_14841# a_643_15213# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2153 a_127_3207# a_7331_4818# a_6485_6328# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X2154 a_127_3207# a_14239_10305# a_14407_10207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2155 a_13281_11571# a_12586_11811# a_13199_11571# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2156 a_12586_327# a_13435_995# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2157 a_14079_13721# div_out2_3 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2158 a_1371_9913# a_11903_7763# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2159 a_6185_3433# a_9585_3209# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X2160 a_1673_9939# a_1507_9939# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2161 a_2442_513# a_2316_415# a_2038_399# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2162 a_12803_14835# a_12854_15379# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2163 w_62_9065# a_2754_9627# a_3250_9395# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X2164 a_10073_4858# a_9097_5098# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.325 ps=1.65 w=1 l=0.15
X2165 a_12183_5294# a_11749_5294# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=0.5
X2166 a_739_15213# a_127_14841# a_643_15213# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2167 a_397_13203# a_534_13383# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2168 w_62_12329# a_12174_11179# a_12179_12115# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2169 w_62_2537# a_12586_1415# a_12528_1601# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X2170 a_12528_14657# a_11989_15353# a_12231_14265# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X2171 a_127_3207# a_15188_396# a_15126_513# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2172 a_13814_10483# a_13375_10489# a_13729_10483# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2173 a_12826_147# a_12498_399# a_12402_299# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2174 a_127_3207# a_2114_2435# a_2072_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2175 w_62_15593# div_out0_3 a_13281_14541# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2176 a_13435_995# a_12854_2323# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2177 a_13435_8611# a_13260_8685# a_13614_8673# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2178 a_3746_11027# a_3660_11179# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2179 a_127_3207# a_12854_10483# a_14125_11937# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2180 a_13743_5587# a_6185_3209# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2181 a_905_15201# a_861_14809# a_739_15213# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2182 a_15126_1601# a_14368_1503# a_14563_1472# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.07245 ps=0.765 w=0.42 l=0.15
X2183 a_127_3207# a_122_923# a_127_697# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2184 a_13260_1069# a_12345_697# a_12913_665# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2185 w_62_15593# a_12586_14471# a_12528_14657# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X2186 a_11279_8265# a_5853_8418# a_11279_7927# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.1125 pd=1.05 as=0.225 ps=2.1 w=0.75 l=0.15
X2187 a_1370_9395# a_127_9401# a_1208_9773# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2188 w_62_2537# enb_0 a_10073_6368# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.65 pd=2.65 as=0.6 ps=4.6 w=2 l=0.15
X2189 a_127_3207# w_62_6889# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2190 a_127_3207# div_out1_3 a_13199_13453# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2191 a_3746_691# a_3617_1387# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2192 a_1317_15213# a_293_14841# a_1208_15213# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2193 a_12913_8281# a_12695_8685# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2194 a_14801_8851# a_12854_9939# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2195 a_127_3207# a_4315_15353# a_3617_14443# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2196 a_631_10091# a_1147_8013# a_1397_8013# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X2197 a_2754_9627# a_2703_8307# a_2880_9761# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2198 a_5377_10189# a_5003_10189# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2199 a_11300_11891# a_11279_12307# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.45 pd=3.6 as=0.225 ps=1.8 w=1.5 l=0.15
X2200 a_548_8673# a_127_7763# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2201 w_62_14505# a_4077_13388# a_5678_14627# w_62_14505# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X2202 a_15188_12633# a_15302_12481# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X2203 a_11658_1235# a_11382_1235# a_11300_1485# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2204 a_14494_513# a_14407_289# a_14090_399# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.0588 ps=0.7 w=0.42 l=0.15
X2205 a_12498_8015# a_12402_9003# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2206 a_3250_12481# a_941_12659# a_3140_12481# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X2207 a_13435_15139# a_13260_15213# a_13614_15201# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2208 a_6185_3209# a_13835_5043# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2054 pd=2.1 as=0.11455 ps=1.08 w=0.79 l=0.15
X2209 a_127_3207# a_2511_1472# a_2442_1601# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2210 a_127_3207# a_14368_415# a_14407_289# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2211 a_3074_9217# a_2355_8993# a_2511_9088# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2212 a_12854_10483# a_12271_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2213 w_62_361# a_12586_327# a_12402_299# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X2214 a_2072_2323# a_1673_2323# a_1946_2689# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2215 a_14806_15067# a_14755_13747# a_14932_15201# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2216 a_127_3207# a_5679_2511# a_5419_2297# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2217 w_62_10153# a_14407_10207# a_14838_10261# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X2218 a_1766_15599# a_2970_15701# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2219 a_15188_11545# a_15302_11393# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2220 a_2245_15155# a_1783_14291# a_397_15531# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X2221 w_62_15593# a_2539_15647# a_2970_15701# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X2222 w_62_13417# a_12913_13721# a_12803_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2223 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=0.59
X2224 a_13435_9699# a_12854_9939# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2225 a_13541_15379# a_13375_15379# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2226 w_62_1449# a_2754_2011# a_3250_1779# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X2227 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2228 a_4533_10189# a_3899_10189# a_4315_9913# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2229 w_62_10153# a_2539_10207# a_2455_10305# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1113 pd=1.37 as=0.0882 ps=0.84 w=0.42 l=0.15
X2230 a_548_11027# a_127_11571# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2231 w_62_361# div_out1_0 a_13281_397# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2232 a_127_3207# w_62_5801# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2233 w_62_6889# a_127_3207# w_62_6889# w_62_6889# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2234 w_62_7977# div_fb1_1 a_1229_8013# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2235 a_127_3207# a_11296_14443# a_11903_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2236 a_12586_7943# a_13435_8611# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2237 a_127_3207# a_13887_8825# a_13835_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X2238 a_127_3207# a_1783_14291# a_2027_14809# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2239 a_13982_15491# a_13814_15745# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2240 a_12265_15531# a_14079_14809# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X2241 w_62_10153# a_3617_11803# a_3981_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2242 a_1225_10715# a_3660_12891# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2243 a_2027_8281# div_fb2_1 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2244 a_127_3207# a_12854_9939# a_12957_9761# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2245 a_12803_14835# a_12345_14841# a_12695_15213# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2246 a_15289_15379# a_15123_15379# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2247 a_947_969# a_403_2573# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2248 a_941_13203# a_350_13355# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2249 a_127_3207# a_1835_7737# a_1783_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X2250 w_62_2537# div_out0_0 a_13281_1485# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2251 a_1370_1779# a_127_1785# a_1208_2157# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2252 a_2442_1601# a_2316_1503# a_2038_1487# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2253 w_62_13417# a_2511_13440# a_2442_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2254 w_62_13417# a_12231_13177# a_12179_13203# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X2255 a_12826_7763# a_12498_8015# a_12402_7915# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2256 a_127_3207# div_fb3_0 a_2245_2099# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2257 a_1147_397# a_534_327# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2258 w_62_1449# a_179_1209# a_127_1235# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X2259 a_1673_2323# a_1507_2323# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2260 a_12854_2323# a_12271_2573# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2261 a_14932_14113# a_13835_13203# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X2262 w_62_10153# a_14732_10189# a_15123_9939# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2263 a_12449_147# a_12586_327# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2264 a_15188_13452# a_15302_13747# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X2265 a_5003_10483# a_2864_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2266 a_127_3207# a_12174_11179# a_12179_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2267 a_14090_1487# a_14407_1377# a_14365_1235# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2268 a_127_3207# a_9097_5098# a_10073_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.325 pd=1.65 as=0.3 ps=2.6 w=1 l=0.15
X2269 w_62_5801# a_127_3207# w_62_5801# w_62_5801# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2270 w_62_15593# a_12271_15629# a_13375_15379# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2271 a_12586_13383# a_13435_14051# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.2087 ps=2.02 w=0.65 l=0.15
X2272 a_12449_13203# a_12586_13383# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2273 a_13814_2689# a_13375_2323# a_13729_2323# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0621 pd=0.705 as=0.0813 ps=0.83 w=0.36 l=0.15
X2274 a_127_3207# a_2754_2011# a_2703_1779# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2275 w_62_2537# a_11749_5294# a_12183_5294# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=0.5
X2276 a_2073_11937# a_2038_11703# a_1835_11545# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2277 a_6185_3209# a_13835_5043# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1352 pd=1.56 as=0.0754 ps=0.81 w=0.52 l=0.15
X2278 a_127_3207# a_14407_10457# a_14838_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.1092 ps=1.36 w=0.42 l=0.15
X2279 a_14465_11277# div_out3_2 w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2280 a_3136_396# a_3250_691# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2281 a_13982_10051# a_13814_10305# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2282 a_2749_8851# a_947_8585# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2283 a_127_3207# a_6185_3209# a_13743_5587# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2284 a_2749_147# a_947_969# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2285 a_127_3207# a_14563_14528# a_14494_14657# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2286 a_739_1069# a_127_697# a_643_1069# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2287 a_774_1235# a_121_2297# a_350_1387# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1092 ps=1.36 w=0.42 l=0.15
X2288 a_15289_2323# a_15123_2323# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2289 w_62_10153# a_14806_11179# a_15302_11393# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X2290 a_12271_15629# a_12499_15531# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.089375 ps=0.925 w=0.65 l=0.15
X2291 a_127_3207# a_13435_2083# a_13369_2157# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2292 a_13435_2083# a_12854_2323# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2293 a_127_3207# a_12595_9913# a_12271_10189# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2294 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2295 w_62_10153# a_13982_10457# a_13909_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.07665 ps=0.785 w=0.42 l=0.15
X2296 w_62_6889# a_127_3207# w_62_6889# w_62_6889# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2297 a_127_3207# a_947_14025# a_905_15201# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2298 w_62_10153# a_11989_9913# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2299 a_1208_15213# a_127_14841# a_861_14809# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2300 w_62_13417# a_534_13383# a_350_13355# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X2301 a_127_3207# a_14806_15067# a_14755_14835# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2302 a_14932_8673# a_13835_7763# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X2303 a_13634_2543# a_14838_2645# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2304 a_2114_10051# a_1946_10305# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2305 a_397_10091# a_2027_9369# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X2306 a_3079_11027# a_2703_12115# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2307 a_127_3207# a_5853_802# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=3.3 pd=22.6 as=0 ps=0 w=11 l=2
X2308 a_1562_15201# a_947_14025# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2309 a_2880_11027# a_1783_11571# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X2310 a_15192_14835# a_13835_14291# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X2311 a_5377_10483# a_5003_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2312 a_179_121# a_350_299# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X2313 a_14563_8000# a_14407_7905# a_14708_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2314 a_2027_665# a_1783_147# a_2413_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2315 a_13940_2323# a_13541_2323# a_13814_2689# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0696 pd=0.765 as=0.0621 ps=0.705 w=0.36 l=0.15
X2316 w_62_10153# a_13435_9699# a_13422_9395# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2317 a_3763_8825# a_5419_9913# a_5377_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2318 a_14324_13569# a_13887_13177# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2319 w_62_361# a_2754_923# a_2703_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2320 w_62_13417# a_3136_13452# a_3074_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2321 a_567_2573# a_535_2475# a_485_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2322 a_10073_7110# a_9567_6368# a_6185_3321# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.325 pd=1.65 as=0.3 ps=2.6 w=1 l=0.5
X2323 a_4825_10189# a_4315_9913# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2324 w_62_9065# a_534_9031# a_350_9003# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X2325 w_62_13417# a_14368_13471# a_14407_13345# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2326 a_2114_15491# a_1946_15745# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.178875 ps=1.26 w=0.75 l=0.15
X2327 a_9193_4818# a_6485_5594# a_8019_4858# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=0.5
X2328 a_15188_9100# a_15302_9395# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X2329 a_3379_10821# a_1225_10715# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2330 a_13729_2323# a_13634_2543# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2331 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2332 a_5853_802# a_3763_1209# a_5678_414# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=0.15
X2333 w_62_11241# a_861_11269# a_751_11393# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.07035 pd=0.755 as=0.1155 ps=0.97 w=0.42 l=0.15
X2334 a_13260_11027# a_12179_11027# a_12913_11269# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2335 a_4533_10483# a_3899_10483# a_4315_10457# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2336 a_13435_12089# a_12854_10483# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2337 a_14239_2689# a_13541_2323# a_13982_2435# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2338 a_2313_14291# a_1835_14265# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2339 a_12435_2573# a_12403_2475# a_12353_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.19 pd=1.38 as=0.13 ps=1.26 w=1 l=0.15
X2340 a_127_3207# w_62_3625# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2341 a_3660_2011# a_3763_1209# a_3709_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2342 a_11296_14443# a_11658_14291# a_11300_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2343 a_6185_3545# a_9585_3321# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X2344 w_62_7977# a_11296_9003# a_11903_7763# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2345 a_2656_9217# a_2442_9217# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2346 w_62_3625# a_127_3207# w_62_3625# w_62_3625# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2347 a_3981_10189# a_3657_9939# a_3899_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2348 a_1946_10305# a_1673_9939# a_1861_9939# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2349 a_11300_14291# a_11279_13705# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.45 pd=3.6 as=0.225 ps=1.8 w=1.5 l=0.15
X2350 a_11279_7927# a_5853_8418# a_11279_8265# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.225 pd=2.1 as=0.1125 ps=1.05 w=0.75 l=0.15
X2351 a_2057_12365# a_1783_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2352 a_3140_11393# a_1783_11571# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X2353 a_2754_13979# a_1783_13203# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.14075 ps=1.325 w=0.42 l=0.15
X2354 a_127_3207# a_947_14025# a_2073_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2355 a_127_3207# a_6422_13265# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.6 pd=4.3 as=0 ps=0 w=4 l=6
X2356 a_127_3207# a_2511_13440# a_2442_13569# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2357 a_2371_15745# a_1673_15379# a_2114_15491# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0684 pd=0.74 as=0.0989 ps=0.995 w=0.36 l=0.15
X2358 a_12993_13203# a_12402_13355# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.14075 ps=1.325 w=1 l=0.15
X2359 w_62_13417# a_941_13203# a_2754_13979# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X2360 a_3660_15067# a_3763_14265# a_3709_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2361 a_1370_14835# a_127_14841# a_1208_15213# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2362 a_2027_12300# a_1783_12659# a_2413_12365# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2363 a_13814_10305# a_13541_9939# a_13729_9939# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.05775 ps=0.695 w=0.42 l=0.15
X2364 a_14365_147# a_13887_121# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2365 a_2245_11027# a_1783_11571# a_397_10715# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X2366 a_127_3207# a_14368_12775# a_14407_12901# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2367 a_3136_8012# a_3250_8307# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X2368 w_62_15593# a_12854_15379# a_13887_14265# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2369 a_12265_2475# a_14079_1753# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X2370 w_62_10153# a_14732_10483# a_15123_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2371 w_62_14505# a_1225_15531# a_4971_13388# w_62_14505# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1 as=0.15 ps=1.6 w=0.5 l=0.15
X2372 w_62_2537# a_13435_2083# a_13422_1779# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2373 a_127_3207# a_12271_15629# a_13375_15379# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2374 a_3379_9967# a_1225_10091# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2375 a_127_3207# a_1783_11571# a_2027_11212# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2376 a_13435_995# a_13260_1069# a_13614_1057# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2377 a_127_3207# a_259_10457# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2378 a_12265_10715# a_14079_11212# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X2379 a_15188_1484# a_15302_1779# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.23605 ps=1.765 w=1 l=0.15
X2380 a_12695_9773# a_12345_9401# a_12600_9761# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2381 a_7331_5294# a_9097_5098# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.15 pd=1.6 as=0.075 ps=0.8 w=0.5 l=0.15
X2382 a_127_3207# a_3136_13452# a_3074_13569# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2205 pd=1.89 as=0.066 ps=0.745 w=0.42 l=0.15
X2383 w_62_12329# a_534_12899# a_350_12891# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X2384 w_62_10153# div_out3_1 a_14109_9395# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2385 a_127_3207# div_out3_3 a_14297_15155# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2386 a_127_3207# div_fb0_3 a_1147_14541# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2387 a_12586_11811# a_13435_11001# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3012 ps=2.66 w=1 l=0.15
X2388 w_62_2537# a_9097_5098# a_11630_6516# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2389 a_127_3207# a_12854_15379# a_12957_15201# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2390 a_12402_13355# a_12498_13455# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X2391 w_62_13417# a_12586_13383# a_12402_13355# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X2392 a_14801_1235# a_12854_2323# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2393 a_2316_14559# a_122_13979# w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2394 a_941_12659# a_350_12891# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2395 a_2754_2011# a_2703_691# a_2880_2145# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2396 a_14079_1753# div_out3_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2397 a_548_1057# a_127_147# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2398 a_1383_11001# a_1208_11027# a_1562_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.06405 ps=0.725 w=0.42 l=0.15
X2399 a_14090_399# a_14407_289# a_14365_147# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2400 a_127_3207# a_12231_12633# a_12179_12659# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2401 a_13909_15745# a_13375_15379# a_13814_15745# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.06825 ps=0.745 w=0.42 l=0.15
X2402 a_14324_12659# a_13887_12633# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2403 a_8019_6368# a_9193_6328# a_9151_7110# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.3 as=0.105 ps=1.21 w=1 l=0.5
X2404 a_14494_13569# a_14368_13471# a_14090_13455# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2405 w_62_12329# a_3136_12633# a_3074_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2406 a_127_3207# a_6422_209# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=1.2 pd=8.6 as=0 ps=0 w=4 l=6
X2407 a_2057_13747# a_1783_13203# w_62_13417# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2408 a_14368_12775# a_12174_11179# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2409 a_2754_11179# a_2703_12115# a_2880_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0441 ps=0.63 w=0.42 l=0.15
X2410 a_3763_11545# a_5419_10457# a_5377_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2411 a_3074_1601# a_2355_1377# a_2511_1472# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2412 a_127_3207# a_7331_4818# a_6485_6328# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X2413 w_62_13417# a_4910_13976# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X2414 a_127_3207# a_11296_9003# a_11903_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0754 pd=0.81 as=0.1352 ps=1.56 w=0.52 l=0.15
X2415 w_62_12329# a_14806_12267# a_14755_12115# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2416 a_861_665# a_643_1069# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.12915 pd=1.185 as=0.2184 ps=2.2 w=0.84 l=0.15
X2417 a_14125_8851# a_14090_9103# a_13887_8825# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2418 a_2272_9217# a_1835_8825# w_62_9065# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2419 a_13887_121# a_14090_399# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2420 a_4825_10483# a_4315_10457# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2421 a_2511_384# a_2316_415# a_2821_147# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2422 a_12600_12115# a_12179_12659# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.2205 ps=1.89 w=0.42 l=0.15
X2423 a_12402_9003# a_11989_9913# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X2424 a_2027_13721# a_1783_13203# a_2413_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2425 a_14708_1601# a_14494_1601# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07035 ps=0.755 w=0.42 l=0.15
X2426 a_4575_10127# a_3746_9395# a_4825_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2427 w_62_11241# a_534_11811# a_350_11803# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X2428 a_739_12115# a_127_12115# a_643_12115# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.1401 pd=1.1 as=0.0594 ps=0.69 w=0.36 l=0.15
X2429 a_2073_7763# a_2038_8015# a_1835_7737# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2430 w_62_1449# a_1835_1209# a_1783_1235# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.3012 pd=2.66 as=0.26 ps=2.52 w=1 l=0.15
X2431 a_2316_9119# a_122_8539# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2432 a_4971_12724# a_4137_12618# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X2433 a_127_3207# a_14806_11179# a_14755_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2434 a_13281_397# a_12586_327# a_13199_397# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2435 a_127_3207# a_13887_1209# a_13835_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X2436 a_12957_14113# a_12913_13721# a_12791_14125# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2437 w_62_13417# a_13435_14051# a_13422_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2438 a_127_3207# w_62_6889# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2439 a_446_12633# a_350_11803# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2440 a_127_3207# w_62_3625# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=4.73
X2441 a_9151_6368# enb_0 w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.21 pd=2.21 as=0.6 ps=4.6 w=2 l=0.15
X2442 a_13449_9101# div_out0_1 w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2443 a_12854_15379# a_12271_15629# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2444 a_1673_10489# a_1507_10489# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2445 a_127_3207# a_12231_11545# a_12179_11571# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2446 a_12600_8673# a_12179_7763# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0651 pd=0.73 as=0.1092 ps=1.36 w=0.42 l=0.15
X2447 a_3981_10483# a_3657_10483# a_3899_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2448 a_14324_11571# a_13887_11545# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2449 a_127_3207# a_12854_2323# a_12957_2145# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0441 ps=0.63 w=0.42 l=0.15
X2450 w_62_11241# a_3136_11545# a_3074_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2451 w_62_2537# div_out3_0 a_14109_1779# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2452 w_62_3625# a_127_3207# w_62_3625# w_62_3625# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2453 a_127_3207# a_13835_8851# a_14079_9369# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2454 a_1317_12115# a_293_12115# a_1208_12115# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2455 w_62_13417# a_12174_13979# a_12179_13753# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2456 a_12913_12357# a_12695_12115# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2457 a_947_11001# a_403_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2458 w_62_361# a_2754_923# a_3250_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X2459 a_5419_10457# a_5003_10483# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2460 w_62_1449# a_122_923# a_127_1785# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2461 w_62_2537# enb_0 a_9887_6368# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.21 ps=2.21 w=2 l=0.15
X2462 a_293_13753# a_127_13753# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2463 a_127_3207# a_3519_10499# a_3465_10821# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1118 pd=1.04 as=0.0567 ps=0.69 w=0.42 l=0.15
X2464 a_1835_1209# a_2038_1487# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1134 ps=1.38 w=0.42 l=0.15
X2465 a_15302_11393# a_14806_11179# a_15131_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2466 a_2455_10483# a_1673_10489# a_2371_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2467 w_62_15593# a_3617_14443# a_3981_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2468 a_14732_10189# a_14407_10207# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2469 a_14368_14559# a_12174_13979# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2470 w_62_15593# a_121_15353# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2471 w_62_4713# a_127_3207# w_62_4713# w_62_4713# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2472 a_127_3207# w_62_5801# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=1.05
X2473 a_2749_1235# a_947_969# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2474 w_62_6889# a_127_3207# w_62_6889# w_62_6889# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2475 a_127_3207# a_534_9031# a_774_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X2476 w_62_13417# a_14806_13979# a_14755_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.26 ps=2.52 w=1 l=0.15
X2477 a_127_3207# w_62_2537# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.143 pd=1.62 as=0 ps=0 w=0.55 l=0.59
X2478 a_127_3207# a_2539_10457# a_2497_10861# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2479 a_403_15629# a_397_15531# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
X2480 a_751_11393# a_947_11001# w_62_11241# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2481 a_127_3207# a_13982_2435# a_13940_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0696 ps=0.765 w=0.42 l=0.15
X2482 a_12402_12891# a_12498_12633# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X2483 a_14323_10483# a_13541_10489# a_14239_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.0567 ps=0.69 w=0.42 l=0.15
X2484 w_62_7977# a_12586_7943# a_12402_7915# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X2485 a_179_1209# a_350_1387# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X2486 w_62_12329# a_12586_12899# a_12402_12891# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X2487 a_127_3207# a_4575_2511# a_4315_2297# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2488 w_62_7977# a_1208_8685# a_1383_8611# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2489 a_127_3207# a_6185_3209# a_13743_5587# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2490 w_62_5801# a_127_3207# w_62_5801# w_62_5801# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2491 a_14932_1057# a_13835_147# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.097 ps=0.975 w=0.42 l=0.15
X2492 a_11382_8851# a_11296_9003# a_11300_9101# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2493 a_2821_13025# a_2442_12659# a_2749_13025# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2494 a_1397_8851# div_fb0_1 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2495 a_127_3207# a_535_10091# a_403_10189# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X2496 a_127_3207# a_5853_11873# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=3.3 pd=22.6 as=0 ps=0 w=11 l=2
X2497 a_1317_2323# a_1225_2475# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2498 a_127_3207# a_14563_8000# a_14494_8129# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1346 pd=1.15 as=0.0999 ps=0.985 w=0.64 l=0.15
X2499 a_3709_14291# a_3617_14443# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2500 a_751_11393# a_293_11027# a_643_11027# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2501 a_13185_9939# a_1225_10091# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2502 w_62_9065# a_947_8585# a_1835_8825# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2503 a_11658_14291# a_11382_14291# a_11300_14541# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.26 ps=2.52 w=1 l=0.15
X2504 a_2057_11277# a_2027_11212# a_397_10715# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X2505 a_14090_13455# a_14407_13345# a_14365_13203# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2506 a_12993_12659# a_12402_12891# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2507 a_14324_1601# a_13887_1209# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0819 ps=0.81 w=0.42 l=0.15
X2508 a_293_697# a_127_697# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2509 w_62_2537# a_12595_2297# a_12541_2573# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2510 a_2413_691# div_fb2_0 w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2511 a_673_10189# a_631_10091# a_567_10189# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X2512 a_6185_3433# a_9585_3657# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
X2513 a_11296_9003# a_11658_8851# a_11300_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2514 w_62_10153# a_12231_8825# a_12179_8851# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X2515 a_127_3207# a_12403_10091# a_12271_10189# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X2516 w_62_12329# div_out2_2 a_14109_12365# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2517 a_12499_2475# a_12586_327# a_13449_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2518 a_127_3207# a_535_15531# a_403_15629# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X2519 w_62_5801# a_127_3207# w_62_5801# w_62_5801# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=1.05
X2520 a_12803_11393# a_12854_10483# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2521 a_15302_12481# a_12993_12659# a_15192_12481# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X2522 a_9151_4858# a_9097_5098# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.105 pd=1.21 as=0.3 ps=2.6 w=1 l=0.15
X2523 a_476_9217# a_121_9913# a_179_8825# w_62_9065# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.0567 ps=0.69 w=0.42 l=0.15
X2524 a_1317_9773# a_293_9401# a_1208_9773# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2525 a_403_10189# a_397_10091# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
X2526 a_12271_10483# a_12265_10715# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
X2527 a_12402_11803# a_11989_10748# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0609 pd=0.71 as=0.1491 ps=1.13 w=0.42 l=0.15
X2528 a_4575_10457# a_3746_11027# a_4825_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2529 a_15188_8012# a_15302_8307# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2530 w_62_10153# a_12586_11811# a_12402_11803# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.14075 pd=1.325 as=0.0609 ps=0.71 w=0.42 l=0.15
X2531 a_2316_1503# a_122_923# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2532 a_127_3207# div_out3_2 a_14297_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2533 a_5377_15629# a_5003_15629# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2534 a_1208_8685# a_127_8313# a_861_8281# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2535 a_12074_7210# a_11654_6816# a_11594_6922# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.15 pd=1.6 as=0.15 ps=1.6 w=0.5 l=2.1
X2536 a_1208_12115# a_293_12115# a_861_12357# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2537 a_127_3207# a_1783_12659# a_3079_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2538 a_14297_15155# a_13835_14291# a_12265_15531# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X2539 a_14090_9103# a_14368_9119# a_14324_9217# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2540 a_1147_14541# a_534_14471# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2541 a_2316_13471# a_122_13979# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2542 a_535_2475# a_2027_665# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.208 ps=1.94 w=0.65 l=0.15
X2543 a_12271_10189# a_12265_10091# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.118625 pd=1.015 as=0.169 ps=1.82 w=0.65 l=0.15
X2544 a_11279_13367# a_5853_13858# a_11279_13705# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.225 pd=2.1 as=0.1125 ps=1.05 w=0.75 l=0.15
X2545 a_12498_12633# a_12402_11803# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2546 a_13260_9773# a_12179_9401# a_12913_9369# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2547 a_14801_147# a_12854_2323# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1346 ps=1.15 w=0.42 l=0.15
X2548 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2549 a_2038_13455# a_2316_13471# a_2272_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2550 a_751_8307# a_947_8585# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2551 a_2245_9715# a_1783_8851# a_397_10091# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X2552 a_127_3207# a_9097_5098# a_9887_4858# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.105 ps=1.21 w=1 l=0.15
X2553 a_13634_15599# a_14838_15701# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2554 a_751_691# a_947_969# w_62_361# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.07035 ps=0.755 w=0.42 l=0.15
X2555 a_2038_8015# a_2316_8031# a_2272_8129# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2556 a_3379_2351# a_1225_2475# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.1176 ps=1.4 w=0.42 l=0.15
X2557 w_62_7977# a_4910_8536# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=1.8
X2558 w_62_15593# a_14407_15647# a_14838_15701# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.1664 ps=1.8 w=0.64 l=0.15
X2559 a_1208_12115# a_127_12115# a_861_12357# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0999 ps=0.985 w=0.36 l=0.15
X2560 a_4533_15629# a_3899_15629# a_4315_15353# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2561 w_62_2537# a_127_3207# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.2262 pd=2.26 as=0 ps=0 w=0.87 l=4.73
X2562 a_127_3207# a_12403_10715# a_12271_10483# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.089375 pd=0.925 as=0.118625 ps=1.015 w=0.65 l=0.15
X2563 a_14494_12659# a_14368_12775# a_14090_12791# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0999 pd=0.985 as=0.0711 ps=0.755 w=0.36 l=0.15
X2564 a_127_3207# a_12231_121# a_12179_147# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2565 a_12231_14265# a_12402_14443# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.23605 ps=1.765 w=0.42 l=0.15
X2566 w_62_2537# enb_0 a_10097_3881# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.45 pd=3.6 as=0.225 ps=1.8 w=1.5 l=0.15
X2567 a_3250_8307# a_941_7763# a_3140_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X2568 w_62_12329# a_1208_12115# a_1383_12089# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.1134 pd=1.38 as=0.0567 ps=0.69 w=0.42 l=0.15
X2569 w_62_13417# a_14563_13440# a_14494_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.2184 pd=2.2 as=0.12915 ps=1.185 w=0.84 l=0.15
X2570 a_10097_3881# enb_0 w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.225 pd=1.8 as=0.45 ps=3.6 w=1.5 l=0.15
X2571 a_14732_10483# a_14407_10457# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2572 w_62_13417# div_out2_3 a_14109_13747# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2573 a_127_3207# a_12271_2573# a_13375_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2574 a_13729_10483# a_13634_10647# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.1092 ps=1.36 w=0.42 l=0.15
X2575 a_446_8015# a_350_9003# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2576 w_62_15593# a_12586_14471# a_13449_14541# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2577 a_12695_2157# a_12345_1785# a_12600_2145# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.066 ps=0.745 w=0.36 l=0.15
X2578 a_3763_8825# a_5003_10189# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2579 w_62_361# a_12586_327# a_12528_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.084 ps=0.82 w=0.42 l=0.15
X2580 a_127_3207# a_121_10748# a_397_11937# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2581 a_5175_12724# a_4971_12724# a_4077_12724# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.075 pd=0.8 as=0.15 ps=1.6 w=0.5 l=0.15
X2582 a_2511_384# a_2355_289# a_2656_513# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.1155 ps=0.97 w=0.42 l=0.15
X2583 a_13281_8013# a_12586_7943# a_13199_8013# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2584 a_14125_11937# a_14090_11703# a_13887_11545# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2585 a_127_3207# a_1835_14265# a_1783_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.2087 pd=2.02 as=0.169 ps=1.82 w=0.65 l=0.15
X2586 w_62_10153# a_403_10483# a_1507_10489# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X2587 w_62_2537# a_12854_2323# a_13887_1209# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.0819 pd=0.81 as=0.0567 ps=0.69 w=0.42 l=0.15
X2588 a_293_8313# a_127_8313# w_62_7977# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X2589 a_3079_9761# a_2703_8307# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2590 a_14873_8851# a_14494_9217# a_14801_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1401 pd=1.1 as=0.0441 ps=0.63 w=0.42 l=0.15
X2591 w_62_15593# a_14732_15629# a_15123_15379# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2592 a_12499_15531# a_12586_13383# a_13449_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2593 a_127_3207# a_727_2297# a_403_2573# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2594 a_127_3207# div_out2_1 a_14297_8627# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2595 a_14365_8851# a_13887_8825# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0669 pd=0.75 as=0.12495 ps=1.015 w=0.42 l=0.15
X2596 a_4137_7908# a_4077_7948# a_4711_9187# w_62_9065# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=1
X2597 a_4137_13348# a_4077_13388# a_4711_14627# w_62_14505# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=1
X2598 a_12803_11393# a_12345_11027# a_12695_11027# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2599 w_62_7977# a_12993_7763# a_14806_8539# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X2600 a_13982_10051# a_13814_10305# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.12095 ps=1.085 w=0.64 l=0.15
X2601 a_12174_11179# a_1371_10457# a_13185_10803# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2602 a_2027_12300# div_fb2_2 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.08775 ps=0.92 w=0.65 l=0.15
X2603 a_127_3207# a_122_13979# a_127_13753# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X2604 a_673_10483# a_631_10715# a_567_10483# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.19 ps=1.38 w=1 l=0.15
X2605 a_14297_2099# a_13835_1235# a_12265_2475# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X2606 a_14732_15629# a_14407_15647# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2607 w_62_361# a_179_121# a_127_147# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.26 ps=2.52 w=1 l=0.15
X2608 a_15131_11027# a_14755_12115# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2609 a_13614_15201# a_12854_15379# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.12495 ps=1.015 w=0.42 l=0.15
X2610 a_9887_5400# a_9193_4818# a_8199_4858# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.21 pd=2.21 as=0.3 ps=2.3 w=2 l=0.5
X2611 a_14125_1235# a_14090_1487# a_13887_1209# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.06405 pd=0.725 as=0.1092 ps=1.36 w=0.42 l=0.15
X2612 w_62_10153# a_14239_10305# a_14407_10207# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.27 ps=2.54 w=1 l=0.15
X2613 a_4315_9913# a_3899_10189# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2614 a_1861_9939# a_1766_10159# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2615 a_14109_9395# a_14079_9369# a_12265_10091# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X2616 a_941_147# a_350_299# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.097 ps=0.975 w=0.65 l=0.15
X2617 w_62_2537# a_7331_5294# a_11654_6816# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.6 ps=4.6 w=2 l=1
X2618 a_12913_13721# a_12695_14125# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0999 pd=0.985 as=0.1346 ps=1.15 w=0.64 l=0.15
X2619 w_62_13417# a_15188_13452# a_15126_13569# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.0651 ps=0.73 w=0.42 l=0.15
X2620 a_12127_15573# a_127_3207# sky130_fd_pr__res_generic_po w=0.48 l=0.045
X2621 a_127_3207# a_4137_7908# a_5678_8030# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.3 ps=2.6 w=1 l=1
X2622 a_127_3207# a_121_9913# a_397_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2623 a_2316_1503# a_122_923# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2624 a_12695_9773# a_12179_9401# a_12600_9761# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.07245 pd=0.765 as=0.0651 ps=0.73 w=0.42 l=0.15
X2625 w_62_10153# a_1371_9913# a_122_8539# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.135 ps=1.27 w=1 l=0.15
X2626 a_9567_6368# a_6185_3321# sky130_fd_pr__cap_mim_m3_1 l=6 w=7
X2627 a_2497_2323# a_1507_2323# a_2371_2689# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2628 a_127_3207# a_13435_15139# a_13369_15213# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2629 a_5225_9261# a_4971_7948# a_4971_7948# w_62_9065# sky130_fd_pr__pfet_01v8 ad=0.125 pd=1 as=0.15 ps=1.6 w=0.5 l=0.15
X2630 a_14365_9939# a_13375_9939# a_14239_10305# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2631 a_2038_12791# a_2316_12775# a_2272_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2632 a_12595_9913# a_12586_9031# a_13449_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.25025 pd=1.42 as=0.08775 ps=0.92 w=0.65 l=0.15
X2633 a_3763_14265# a_5419_15353# a_5377_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.105 ps=1.21 w=1 l=0.15
X2634 a_3074_11571# a_2355_11813# a_2511_11545# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0594 ps=0.69 w=0.36 l=0.15
X2635 a_13260_15213# a_12345_14841# a_12913_14809# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.12915 ps=1.185 w=0.42 l=0.15
X2636 a_15302_8307# a_14806_8539# a_15131_8673# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X2637 a_4825_15629# a_4315_15353# w_62_15593# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2638 a_127_3207# a_12586_7943# a_12826_7763# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X2639 a_14090_12791# a_14407_12901# a_14365_13025# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0711 pd=0.755 as=0.0669 ps=0.75 w=0.36 l=0.15
X2640 w_62_12329# div_out1_2 a_13281_12659# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2641 a_5419_2297# a_5003_2573# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X2642 a_127_3207# a_2539_2591# a_2497_2323# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2643 a_2413_14835# div_fb3_3 w_62_14505# w_62_14505# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2644 a_14109_12365# a_13835_12659# w_62_12329# w_62_12329# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2645 a_127_3207# a_12498_13455# a_12449_13203# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.0567 ps=0.69 w=0.42 l=0.15
X2646 a_127_3207# a_14407_10207# a_14365_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.066 ps=0.745 w=0.42 l=0.15
X2647 a_15192_11393# a_13835_11571# w_62_10153# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.084 pd=0.82 as=0.1491 ps=1.13 w=0.42 l=0.15
X2648 a_4137_12618# a_4137_12618# a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.3 pd=2.6 as=0.15 ps=1.3 w=1 l=1
X2649 a_13743_5587# a_6185_3209# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2650 a_127_3207# a_947_8585# a_2073_8851# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2651 a_127_3207# a_12854_15379# a_14125_14291# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.06405 ps=0.725 w=0.42 l=0.15
X2652 a_3660_2011# a_3617_1387# w_62_1449# w_62_1449# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X2653 a_2511_11545# a_2316_11687# a_2821_11937# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0594 pd=0.69 as=0.1401 ps=1.1 w=0.36 l=0.15
X2654 a_13369_14125# a_12345_13753# a_13260_14125# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.0669 pd=0.75 as=0.0711 ps=0.755 w=0.36 l=0.15
X2655 a_2497_15379# a_1507_15379# a_2371_15745# a_127_3207# sky130_fd_pr__special_nfet_01v8 ad=0.066 pd=0.745 as=0.0684 ps=0.74 w=0.36 l=0.15
X2656 a_3250_691# a_941_147# a_3140_691# w_62_361# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.084 ps=0.82 w=0.42 l=0.15
X2657 w_62_10153# a_15123_9939# a_15289_9939# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.135 ps=1.27 w=1 l=0.15
X2658 a_12803_9395# a_12345_9401# a_12695_9773# w_62_10153# sky130_fd_pr__pfet_01v8_hvt ad=0.1155 pd=0.97 as=0.07245 ps=0.765 w=0.42 l=0.15
X2659 w_62_2537# a_12183_5294# a_11749_5294# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.3 pd=2.3 as=0.6 ps=4.6 w=2 l=0.5
X2660 a_127_3207# a_3746_14835# a_5679_15567# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2661 a_3981_15629# a_3657_15379# a_3899_15629# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.105 pd=1.21 as=0.26 ps=2.52 w=1 l=0.15
X2662 a_127_3207# a_1383_12089# a_1317_12115# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.12495 pd=1.015 as=0.0669 ps=0.75 w=0.42 l=0.15
X2663 a_13422_14835# a_12179_14841# a_13260_15213# w_62_15593# sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0588 ps=0.7 w=0.42 l=0.15
X2664 a_14297_11027# a_13835_11571# a_12265_10715# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.25025 ps=1.42 w=0.65 l=0.15
X2665 a_2038_11703# a_2316_11687# a_2272_11571# w_62_11241# sky130_fd_pr__pfet_01v8_hvt ad=0.0588 pd=0.7 as=0.0567 ps=0.69 w=0.42 l=0.15
X2666 w_62_13417# a_11296_14443# a_11903_13203# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.11455 pd=1.08 as=0.2054 ps=2.1 w=0.79 l=0.15
X2667 a_127_3207# a_534_1415# a_774_1235# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.0441 ps=0.63 w=0.42 l=0.15
X2668 a_11279_12307# a_5853_11873# a_11279_10695# a_127_3207# sky130_fd_pr__nfet_01v8_lvt ad=0.1125 pd=1.05 as=0.225 ps=2.1 w=0.75 l=0.15
X2669 a_127_3207# a_14806_9627# a_14755_9395# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X2670 a_12499_15531# a_13199_13453# a_13449_13453# w_62_13417# sky130_fd_pr__pfet_01v8_hvt ad=0.3 pd=2.6 as=0.26 ps=2.52 w=1 l=0.15
X2671 a_9097_5098# enb_0 a_127_3207# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.169 ps=1.82 w=0.65 l=0.15
X2672 w_62_7977# a_14806_8539# a_15302_8307# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.23605 pd=1.765 as=0.0567 ps=0.69 w=0.42 l=0.15
X2673 a_14109_1779# a_14079_1753# a_12265_2475# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.26 pd=2.52 as=0.3 ps=2.6 w=1 l=0.15
X2674 a_11749_5294# a_11749_5294# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8 ad=0.6 pd=4.6 as=0.3 ps=2.3 w=2 l=0.5
X2675 a_127_3207# a_15123_9939# a_15289_9939# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X2676 w_62_7977# a_941_7763# a_2754_8539# w_62_7977# sky130_fd_pr__pfet_01v8_hvt ad=0.1491 pd=1.13 as=0.0609 ps=0.71 w=0.42 l=0.15
X2677 a_13729_2323# a_13634_2543# w_62_2537# w_62_2537# sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.1092 ps=1.36 w=0.42 l=0.15
X2678 a_905_11027# a_861_11269# a_739_11027# a_127_3207# sky130_fd_pr__nfet_01v8 ad=0.0441 pd=0.63 as=0.1401 ps=1.1 w=0.42 l=0.15
X2679 a_6185_3545# a_9585_3769# a_127_3207# sky130_fd_pr__res_xhigh_po_0p35 l=15
.ends

.subckt tt_um_tiny_pll VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4]
+ uo_out[5] uo_out[6] uo_out[7]
Xsky130_fd_sc_hd__decap_6_46 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_24 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_35 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkbuf_1_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__clkbuf_1_7/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_3_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__clkbuf_2_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_3/A sky130_fd_sc_hd__mux2_1_4/A1
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__dfrtp_1_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_10/A sky130_fd_sc_hd__mux2_1_33/X
+ sky130_fd_sc_hd__clkbuf_2_8/A sky130_fd_sc_hd__mux4_2_0/S0 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfrtp_1_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_4/X sky130_fd_sc_hd__mux2_1_21/X
+ sky130_fd_sc_hd__clkbuf_2_5/X tt08_integration_0/div_fb2_2 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_209 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_1_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_4/X sky130_fd_sc_hd__mux2_1_4/A1
+ sky130_fd_sc_hd__mux2_1_5/S sky130_fd_sc_hd__mux2_1_4/A0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_6_47 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_36 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkbuf_1_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_0/A sky130_fd_sc_hd__clkbuf_2_7/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_3_26 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__clkbuf_2_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__nand4b_1_0/B sky130_fd_sc_hd__nor4b_4_1/C
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__dfrtp_1_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__dfstp_1_10/CLK sky130_fd_sc_hd__mux2_1_37/X
+ sky130_fd_sc_hd__clkbuf_2_6/X sky130_fd_sc_hd__mux4_2_3/S1 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfrtp_1_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_6/X sky130_fd_sc_hd__mux2_1_17/X
+ sky130_fd_sc_hd__clkbuf_2_5/A tt08_integration_0/div_fb3_2 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__mux2_1_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_5/X sky130_fd_sc_hd__buf_2_6/X
+ sky130_fd_sc_hd__mux2_1_5/S sky130_fd_sc_hd__mux2_1_5/A0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_6_48 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_26 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkbuf_1_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__clkbuf_1_9/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_3_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_16 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_ef_sc_hd__decap_12_190 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_1_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__dfstp_1_10/CLK sky130_fd_sc_hd__mux2_1_36/X
+ sky130_fd_sc_hd__clkbuf_2_7/A tt08_integration_0/div_out3_3 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfrtp_1_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_4/X sky130_fd_sc_hd__mux2_1_16/X
+ sky130_fd_sc_hd__clkbuf_2_5/X tt08_integration_0/div_fb1_2 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__nand4b_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_31/S sky130_fd_sc_hd__nor4bb_1_0/A
+ sky130_fd_sc_hd__nand4b_1_0/B sky130_fd_sc_hd__buf_2_9/A sky130_fd_sc_hd__buf_2_8/A
+ sky130_fd_sc_hd__nand4b_1
Xsky130_fd_sc_hd__dfstp_1_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__mux2_1_5/A0 sky130_fd_sc_hd__clkbuf_2_0/X
+ sky130_fd_sc_hd__mux2_1_5/X sky130_fd_sc_hd__clkbuf_1_0/X sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__mux2_1_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_6/X sky130_fd_sc_hd__buf_2_1/X
+ sky130_fd_sc_hd__nor4_4_0/Y tt08_integration_0/div_fb1_0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_6_49 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_16 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_ef_sc_hd__decap_12_350 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_28 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_ef_sc_hd__decap_12_180 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_191 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_1_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__dfstp_1_10/CLK sky130_fd_sc_hd__mux2_1_39/X
+ sky130_fd_sc_hd__clkbuf_2_6/X tt08_integration_0/div_out1_3 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfrtp_1_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__mux2_1_19/X
+ sky130_fd_sc_hd__clkbuf_2_2/X tt08_integration_0/div_fb1_3 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfstp_1_1 VPWR VGND VGND VPWR tt08_integration_0/enb_0 sky130_fd_sc_hd__clkbuf_2_0/X
+ sky130_fd_sc_hd__mux2_1_2/X sky130_fd_sc_hd__clkbuf_1_0/X sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__mux2_1_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_7/X sky130_fd_sc_hd__buf_2_2/X
+ sky130_fd_sc_hd__nor4_4_0/Y tt08_integration_0/div_fb0_0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_6_28 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__dfrtp_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_0/X sky130_fd_sc_hd__mux2_1_1/X
+ sky130_fd_sc_hd__clkbuf_2_0/X sky130_fd_sc_hd__mux2_1_1/A0 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_340 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_ef_sc_hd__decap_12_181 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_170 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_192 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_50 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtp_1_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_10/A sky130_fd_sc_hd__mux2_1_38/X
+ sky130_fd_sc_hd__clkbuf_2_6/X tt08_integration_0/div_out2_3 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfrtp_1_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__dfstp_1_9/CLK sky130_fd_sc_hd__mux2_1_29/X
+ sky130_fd_sc_hd__clkbuf_2_8/X tt08_integration_0/div_out3_2 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfstp_1_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__dfstp_1_2/Q sky130_fd_sc_hd__dfstp_1_2/SET_B
+ sky130_fd_sc_hd__mux2_1_11/X sky130_fd_sc_hd__clkbuf_1_5/X sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__mux2_1_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_8/X sky130_fd_sc_hd__mux2_1_8/A1
+ sky130_fd_sc_hd__mux2_1_9/S tt08_integration_0/div_fb2_1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_6_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__dfrtp_1_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_0/X sky130_fd_sc_hd__mux2_1_0/X
+ sky130_fd_sc_hd__clkbuf_2_0/X sky130_fd_sc_hd__mux2_1_0/A0 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfstp_1_10 VPWR VGND VGND VPWR tt08_integration_0/div_out0_3 sky130_fd_sc_hd__clkbuf_2_6/X
+ sky130_fd_sc_hd__mux2_1_34/X sky130_fd_sc_hd__dfstp_1_10/CLK sky130_fd_sc_hd__dfstp_1
Xsky130_ef_sc_hd__decap_12_330 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_341 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_3_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_ef_sc_hd__decap_12_171 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_160 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_182 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_193 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_51 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtp_1_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__dfstp_1_10/CLK sky130_fd_sc_hd__mux2_1_35/X
+ sky130_fd_sc_hd__clkbuf_2_6/X sky130_fd_sc_hd__mux4_2_3/S0 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfrtp_1_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__mux2_1_25/X
+ sky130_fd_sc_hd__dfstp_1_11/SET_B tt08_integration_0/div_out3_1 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfstp_1_3 VPWR VGND VGND VPWR tt08_integration_0/div_fb0_0 sky130_fd_sc_hd__clkbuf_2_1/X
+ sky130_fd_sc_hd__mux2_1_7/X sky130_fd_sc_hd__dfstp_1_7/CLK sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__mux2_1_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_9/X sky130_fd_sc_hd__buf_2_1/X
+ sky130_fd_sc_hd__mux2_1_9/S tt08_integration_0/div_fb1_1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_6_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__dfrtp_1_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__mux2_1_3/X
+ sky130_fd_sc_hd__dfstp_1_11/SET_B sky130_fd_sc_hd__mux2_1_3/A0 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfstp_1_11 VPWR VGND VGND VPWR tt08_integration_0/div_out0_1 sky130_fd_sc_hd__dfstp_1_11/SET_B
+ sky130_fd_sc_hd__mux2_1_24/X sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__dfstp_1
Xsky130_ef_sc_hd__decap_12_331 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_342 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_320 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4_2/X sky130_fd_sc_hd__mux4_2_3/A0
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_ef_sc_hd__decap_12_183 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_150 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_194 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_161 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_172 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__nor4bb_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_29/S sky130_fd_sc_hd__nor4b_4_1/C
+ sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nor4b_4_0/A sky130_fd_sc_hd__buf_2_8/X
+ sky130_fd_sc_hd__nor4bb_2
Xsky130_fd_sc_hd__decap_4_52 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtp_1_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_5/X sky130_fd_sc_hd__mux2_1_40/X
+ sky130_fd_sc_hd__dfstp_1_2/SET_B tt08_integration_0/div_fb3_1 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfrtp_1_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__dfstp_1_9/CLK sky130_fd_sc_hd__mux2_1_28/X
+ sky130_fd_sc_hd__clkbuf_2_8/X tt08_integration_0/div_out1_2 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfstp_1_4 VPWR VGND VGND VPWR tt08_integration_0/div_fb0_3 sky130_fd_sc_hd__clkbuf_2_2/X
+ sky130_fd_sc_hd__mux2_1_23/X sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__dfrtp_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_0/X sky130_fd_sc_hd__mux2_1_4/X
+ sky130_fd_sc_hd__clkbuf_2_0/X sky130_fd_sc_hd__mux2_1_4/A0 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_332 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_343 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_310 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_321 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_4_2/X sky130_fd_sc_hd__mux4_2_2/A0
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_ef_sc_hd__decap_12_140 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_195 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_184 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_162 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_173 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_151 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_53 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__dfrtp_1_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__dfstp_1_9/CLK sky130_fd_sc_hd__mux2_1_26/X
+ sky130_fd_sc_hd__clkbuf_2_8/X tt08_integration_0/div_out2_2 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfstp_1_5 VPWR VGND VGND VPWR tt08_integration_0/div_fb0_2 sky130_fd_sc_hd__clkbuf_2_5/X
+ sky130_fd_sc_hd__mux2_1_22/X sky130_fd_sc_hd__clkbuf_1_4/X sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__dfrtp_1_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_9/X sky130_fd_sc_hd__mux2_1_41/X
+ sky130_fd_sc_hd__dfstp_1_11/SET_B sky130_fd_sc_hd__dfrtp_1_4/Q sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_333 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_300 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_344 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_311 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_322 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_4_2 VGND VPWR VGND VPWR clk sky130_fd_sc_hd__clkbuf_4_2/X
+ sky130_fd_sc_hd__clkbuf_4
Xsky130_ef_sc_hd__decap_12_130 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_141 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_196 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_174 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_185 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_163 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_152 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_54 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfstp_1_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__dfstp_1_6/Q sky130_fd_sc_hd__clkbuf_2_5/X
+ sky130_fd_sc_hd__mux2_1_13/X sky130_fd_sc_hd__clkbuf_1_4/X sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__dfrtp_1_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_5/X sky130_fd_sc_hd__mux2_1_9/X
+ sky130_fd_sc_hd__dfstp_1_2/SET_B tt08_integration_0/div_fb1_1 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_301 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_312 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_334 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_345 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_323 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_120 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_131 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_142 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_153 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_197 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_186 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_175 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_164 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_0/A sky130_fd_sc_hd__clkbuf_2_0/X
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__decap_4_55 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_44 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfstp_1_7 VPWR VGND VGND VPWR tt08_integration_0/div_fb0_1 sky130_fd_sc_hd__clkbuf_2_1/X
+ sky130_fd_sc_hd__mux2_1_15/X sky130_fd_sc_hd__dfstp_1_7/CLK sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__buf_4_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_0/A uio_oe[5]
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dfrtp_1_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__dfstp_1_7/CLK sky130_fd_sc_hd__mux2_1_10/X
+ sky130_fd_sc_hd__clkbuf_2_1/X tt08_integration_0/div_fb3_0 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_335 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_324 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_302 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_313 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_346 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_110 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_132 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_121 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_165 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_176 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_187 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_154 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_143 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_198 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_2_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_1/A sky130_fd_sc_hd__clkbuf_2_1/X
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__decap_4_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_56 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_45 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfstp_1_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__dfstp_1_8/Q sky130_fd_sc_hd__clkbuf_2_5/X
+ sky130_fd_sc_hd__mux2_1_14/X sky130_fd_sc_hd__clkbuf_1_4/X sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__buf_4_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_1/A uio_oe[6]
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__dfrtp_1_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__dfstp_1_7/CLK sky130_fd_sc_hd__mux2_1_6/X
+ sky130_fd_sc_hd__clkbuf_2_1/X tt08_integration_0/div_fb1_0 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_336 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_303 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_325 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_347 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_314 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_4_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_20/A uo_out[1]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_133 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_100 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_111 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_199 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_122 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_177 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_166 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_155 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_188 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_144 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_2_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_2/A sky130_fd_sc_hd__clkbuf_2_2/X
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__decap_4_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_46 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__dfstp_1_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__dfstp_1_9/Q sky130_fd_sc_hd__clkbuf_2_8/X
+ sky130_fd_sc_hd__mux2_1_27/X sky130_fd_sc_hd__dfstp_1_9/CLK sky130_fd_sc_hd__dfstp_1
Xsky130_fd_sc_hd__buf_4_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_2/A uio_oe[7]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_90 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_1_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__dfstp_1_7/CLK sky130_fd_sc_hd__mux2_1_12/X
+ sky130_fd_sc_hd__clkbuf_2_1/X tt08_integration_0/div_fb2_0 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_304 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_337 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_326 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_348 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_315 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_4_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_10/A uio_out[7]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_0 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_4_21 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_21/A uo_out[5]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_101 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_134 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_123 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_112 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_189 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_167 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_178 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_156 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_145 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_3/A sky130_fd_sc_hd__mux2_1_40/A1
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__decap_4_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_47 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__buf_4_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_3/A uio_oe[4]
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_2_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_0/A
+ sky130_fd_sc_hd__buf_2
Xsky130_ef_sc_hd__decap_12_80 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_91 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__dfrtp_1_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_5/X sky130_fd_sc_hd__mux2_1_8/X
+ sky130_fd_sc_hd__dfstp_1_2/SET_B tt08_integration_0/div_fb2_1 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dlymetal6s2s_1_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__dlymetal6s2s_1_7/A
+ sky130_fd_sc_hd__clkbuf_1_21/X sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_ef_sc_hd__decap_12_338 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_327 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_349 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_316 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_305 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_4_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_11/A uio_out[1]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_1 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_113 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_135 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_124 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_102 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_179 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_168 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_157 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_146 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__and4bb_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__buf_2_0/X
+ sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__mux2_1_43/S
+ sky130_fd_sc_hd__and4bb_1
Xsky130_fd_sc_hd__clkbuf_2_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_9/A sky130_fd_sc_hd__mux2_1_8/A1
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__decap_4_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_48 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__buf_4_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_4/A uo_out[6]
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_2_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_1/X sky130_fd_sc_hd__buf_2_7/A
+ sky130_fd_sc_hd__buf_2
Xsky130_ef_sc_hd__decap_12_92 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_81 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_70 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__dlymetal6s2s_1_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_2/A
+ ui_in[0] sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_fd_sc_hd__mux2_1_40 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_40/X sky130_fd_sc_hd__mux2_1_40/A1
+ sky130_fd_sc_hd__mux2_1_9/S tt08_integration_0/div_fb3_1 sky130_fd_sc_hd__mux2_1
Xsky130_ef_sc_hd__decap_12_317 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_306 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_328 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_339 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_4_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_12/A uio_oe[1]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_2 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_114 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_125 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_136 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_103 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_158 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_169 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_147 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__and4bb_1_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__buf_2_4/X
+ sky130_fd_sc_hd__buf_2_0/X sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__mux2_1_23/S
+ sky130_fd_sc_hd__and4bb_1
Xsky130_fd_sc_hd__clkbuf_2_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_5/A sky130_fd_sc_hd__clkbuf_2_5/X
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__decap_4_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_49 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__buf_4_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_5/A uio_oe[2]
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_2_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_2/X sky130_fd_sc_hd__buf_2_2/A
+ sky130_fd_sc_hd__buf_2
Xsky130_ef_sc_hd__decap_12_82 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_93 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_71 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_60 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__dlymetal6s2s_1_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_8/A
+ sky130_fd_sc_hd__buf_2_0/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_fd_sc_hd__mux2_1_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_30/X sky130_fd_sc_hd__mux4_2_1/S0
+ sky130_fd_sc_hd__mux2_1_31/S sky130_fd_sc_hd__mux2_1_35/A1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_41 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_41/X sky130_fd_sc_hd__buf_2_7/X
+ sky130_fd_sc_hd__mux2_1_3/S sky130_fd_sc_hd__dfrtp_1_4/Q sky130_fd_sc_hd__mux2_1
Xsky130_ef_sc_hd__decap_12_329 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_318 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_307 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_3 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_4_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_13/A uio_out[3]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_115 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_104 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_137 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_126 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_148 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_159 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__and4bb_1_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__nor4b_4_1/C
+ sky130_fd_sc_hd__nor4b_4_0/A sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__mux2_1_3/S
+ sky130_fd_sc_hd__and4bb_1
Xsky130_fd_sc_hd__clkbuf_2_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_8/X sky130_fd_sc_hd__clkbuf_2_6/X
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__decap_4_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__buf_4_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_6/A uio_out[2]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_61 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_50 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_3/X sky130_fd_sc_hd__buf_2_3/A
+ sky130_fd_sc_hd__buf_2
Xsky130_ef_sc_hd__decap_12_94 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_83 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_72 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__dlymetal6s2s_1_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_9/A
+ sky130_fd_sc_hd__buf_2_3/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_fd_sc_hd__mux2_1_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_31/X sky130_fd_sc_hd__mux4_2_1/S1
+ sky130_fd_sc_hd__mux2_1_31/S sky130_fd_sc_hd__mux2_1_37/A1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_42 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_42/X sky130_fd_sc_hd__buf_2_1/X
+ sky130_fd_sc_hd__mux2_1_43/S sky130_fd_sc_hd__mux4_2_2/S1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_20/X sky130_fd_sc_hd__mux2_1_40/A1
+ sky130_fd_sc_hd__mux2_1_23/S tt08_integration_0/div_fb3_3 sky130_fd_sc_hd__mux2_1
Xsky130_ef_sc_hd__decap_12_319 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_308 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_4 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_4_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_14/A uio_out[4]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_105 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_138 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_127 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_116 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_149 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__and4bb_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_9/A sky130_fd_sc_hd__buf_2_8/A
+ sky130_fd_sc_hd__nand4b_1_0/B sky130_fd_sc_hd__nor4bb_1_0/A sky130_fd_sc_hd__mux2_1_33/S
+ sky130_fd_sc_hd__and4bb_1
Xsky130_fd_sc_hd__clkbuf_2_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_7/A sky130_fd_sc_hd__clkbuf_2_8/A
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__decap_4_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_4_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__buf_4_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_7/A uio_out[6]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_84 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_73 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_40 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_95 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_51 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_62 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__buf_2_4/A
+ sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__dlymetal6s2s_1_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_2_7/A
+ sky130_fd_sc_hd__dlymetal6s2s_1_7/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_fd_sc_hd__mux2_1_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_10/X sky130_fd_sc_hd__mux2_1_40/A1
+ sky130_fd_sc_hd__nor4_4_0/Y tt08_integration_0/div_fb3_0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_32 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_32/X sky130_fd_sc_hd__buf_2_7/X
+ sky130_fd_sc_hd__mux2_1_33/S sky130_fd_sc_hd__mux4_2_0/S1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_43 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_43/X sky130_fd_sc_hd__buf_2_2/X
+ sky130_fd_sc_hd__mux2_1_43/S sky130_fd_sc_hd__mux4_2_2/S0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_21/X sky130_fd_sc_hd__mux2_1_8/A1
+ sky130_fd_sc_hd__nor4b_2_0/Y tt08_integration_0/div_fb2_2 sky130_fd_sc_hd__mux2_1
Xsky130_ef_sc_hd__decap_12_309 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_4_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_15/A uio_out[5]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_5 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_3/A ui_in[5]
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_ef_sc_hd__decap_12_117 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_106 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_128 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_139 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_2_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_8/A sky130_fd_sc_hd__clkbuf_2_8/X
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__decap_4_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__decap_3_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__buf_4_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_8/A uo_out[7]
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__buf_2_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__buf_2_5/A
+ sky130_fd_sc_hd__buf_2
Xsky130_ef_sc_hd__decap_12_96 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_85 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_30 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_41 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_74 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_63 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_52 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__dlymetal6s2s_1_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__nand4b_1_0/B
+ sky130_fd_sc_hd__buf_2_4/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_fd_sc_hd__mux2_1_33 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_33/X sky130_fd_sc_hd__buf_2_6/X
+ sky130_fd_sc_hd__mux2_1_33/S sky130_fd_sc_hd__mux4_2_0/S0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_11/X sky130_fd_sc_hd__buf_2_1/X
+ sky130_fd_sc_hd__mux2_1_2/S sky130_fd_sc_hd__dfstp_1_2/Q sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_22/X sky130_fd_sc_hd__buf_2_2/X
+ sky130_fd_sc_hd__nor4b_2_0/Y tt08_integration_0/div_fb0_2 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__buf_4_16 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_16/A uio_oe[3]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_6 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_21/X rst_n
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__clkbuf_1_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_9/A sky130_fd_sc_hd__clkbuf_1_10/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__conb_1_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_8/A sky130_fd_sc_hd__conb_1_10/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_ef_sc_hd__decap_12_118 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_129 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_107 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_2_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_9/A sky130_fd_sc_hd__mux2_1_3/A1
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_ef_sc_hd__decap_12_290 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__buf_4_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_9/A uio_out[0]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_20 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__buf_2_6/A
+ sky130_fd_sc_hd__buf_2
Xsky130_ef_sc_hd__decap_12_31 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_42 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_86 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_75 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_97 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_64 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_53 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_1_23 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_23/X sky130_fd_sc_hd__buf_2_2/X
+ sky130_fd_sc_hd__mux2_1_23/S tt08_integration_0/div_fb0_3 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_34 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_34/X tt08_integration_0/div_out0_3
+ sky130_fd_sc_hd__mux2_1_39/S sky130_fd_sc_hd__buf_2_6/X sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_12/X sky130_fd_sc_hd__mux2_1_8/A1
+ sky130_fd_sc_hd__nor4_4_0/Y tt08_integration_0/div_fb2_0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__nand4b_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__nor4b_4_1/C sky130_fd_sc_hd__mux2_1_39/S
+ sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nor4b_4_0/A
+ sky130_fd_sc_hd__nand4b_2
Xsky130_fd_sc_hd__buf_4_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_17/A uo_out[3]
+ sky130_fd_sc_hd__buf_4
Xsky130_ef_sc_hd__decap_12_7 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__clkbuf_1_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_11/X sky130_fd_sc_hd__clkbuf_1_16/X
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__conb_1_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_7/A sky130_fd_sc_hd__conb_1_11/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_ef_sc_hd__decap_12_119 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_108 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_30 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_ef_sc_hd__decap_12_280 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_291 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_ef_sc_hd__decap_12_10 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_32 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_21 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_43 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__buf_2_7/A
+ sky130_fd_sc_hd__buf_2
Xsky130_ef_sc_hd__decap_12_98 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_87 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_76 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_65 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_54 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_1_35 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_35/X sky130_fd_sc_hd__mux2_1_35/A1
+ sky130_fd_sc_hd__mux2_1_37/S sky130_fd_sc_hd__mux4_2_3/S0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_24 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_24/X sky130_fd_sc_hd__buf_2_6/X
+ sky130_fd_sc_hd__mux2_1_3/S tt08_integration_0/div_out0_1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_13/X sky130_fd_sc_hd__mux2_1_40/A1
+ sky130_fd_sc_hd__mux2_1_2/S sky130_fd_sc_hd__dfstp_1_6/Q sky130_fd_sc_hd__mux2_1
Xsky130_ef_sc_hd__decap_12_8 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_4_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_18/A uo_out[0]
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkbuf_1_12 VGND VPWR VGND VPWR uo_out[4] sky130_fd_sc_hd__clkbuf_1_12/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__conb_1_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_9/A sky130_fd_sc_hd__conb_1_12/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_ef_sc_hd__decap_12_109 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_31 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nor4b_4_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nor4b_4_1/C
+ sky130_fd_sc_hd__nor4b_4_0/A sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__mux2_1_2/S
+ sky130_fd_sc_hd__nor4b_4
Xsky130_ef_sc_hd__decap_12_292 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_270 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_281 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_ef_sc_hd__decap_12_11 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_77 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_33 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_22 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_55 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_66 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_44 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__buf_2_8/A
+ sky130_fd_sc_hd__buf_2
Xsky130_ef_sc_hd__decap_12_99 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_88 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_1_36 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_36/X tt08_integration_0/div_out3_3
+ sky130_fd_sc_hd__mux2_1_39/S sky130_fd_sc_hd__mux2_1_4/A1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_25 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_25/X sky130_fd_sc_hd__mux2_1_4/A1
+ sky130_fd_sc_hd__mux2_1_3/S tt08_integration_0/div_out3_1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_14/X sky130_fd_sc_hd__mux2_1_8/A1
+ sky130_fd_sc_hd__mux2_1_2/S sky130_fd_sc_hd__dfstp_1_8/Q sky130_fd_sc_hd__mux2_1
Xsky130_ef_sc_hd__decap_12_9 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_4_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_4_19/A uo_out[2]
+ sky130_fd_sc_hd__buf_4
Xsky130_fd_sc_hd__clkbuf_1_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_6/A sky130_fd_sc_hd__buf_2_2/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__conb_1_13 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_21/A sky130_fd_sc_hd__conb_1_13/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_21 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__nor4b_4_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_8/X sky130_fd_sc_hd__nor4b_4_0/A
+ sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__nor4b_4_1/C sky130_fd_sc_hd__mux2_1_5/S
+ sky130_fd_sc_hd__nor4b_4
Xsky130_ef_sc_hd__decap_12_293 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_271 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_282 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_260 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_6_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_ef_sc_hd__decap_12_78 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_12 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_23 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_89 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_34 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_56 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_67 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_45 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_9/X sky130_fd_sc_hd__buf_2_9/A
+ sky130_fd_sc_hd__buf_2
Xsky130_fd_sc_hd__mux2_1_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_15/X sky130_fd_sc_hd__buf_2_2/X
+ sky130_fd_sc_hd__mux2_1_9/S tt08_integration_0/div_fb0_1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_26 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_26/X sky130_fd_sc_hd__mux2_1_3/A1
+ sky130_fd_sc_hd__mux2_1_29/S tt08_integration_0/div_out2_2 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_37 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_37/X sky130_fd_sc_hd__mux2_1_37/A1
+ sky130_fd_sc_hd__mux2_1_37/S sky130_fd_sc_hd__mux4_2_3/S1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__clkbuf_1_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_10/A ui_in[1]
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__conb_1_14 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_4/A sky130_fd_sc_hd__conb_1_14/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_33 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_ef_sc_hd__decap_12_283 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_272 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_261 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_250 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_294 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_6_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_ef_sc_hd__decap_12_35 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_24 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_79 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_13 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_46 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_57 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_68 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_1_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_16/X sky130_fd_sc_hd__buf_2_1/X
+ sky130_fd_sc_hd__nor4b_2_0/Y tt08_integration_0/div_fb1_2 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_27 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_27/X sky130_fd_sc_hd__mux2_1_35/A1
+ sky130_fd_sc_hd__mux2_1_29/S sky130_fd_sc_hd__dfstp_1_9/Q sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_38 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_38/X tt08_integration_0/div_out2_3
+ sky130_fd_sc_hd__mux2_1_39/S sky130_fd_sc_hd__mux2_1_3/A1 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__clkbuf_1_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_0/A ui_in[6]
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__conb_1_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_5/A sky130_fd_sc_hd__conb_1_15/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__dlymetal6s2s_1_0 VPWR VGND VGND VPWR sky130_fd_sc_hd__dfstp_1_7/CLK
+ sky130_fd_sc_hd__clkbuf_1_5/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_fd_sc_hd__nor4b_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__buf_2_3/X
+ sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__nor4b_2_0/Y sky130_fd_sc_hd__buf_2_0/X
+ sky130_fd_sc_hd__nor4b_2
Xsky130_ef_sc_hd__decap_12_251 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_262 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_240 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__buf_2_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__buf_2_7/A sky130_fd_sc_hd__buf_2_10/A
+ sky130_fd_sc_hd__buf_2
Xsky130_ef_sc_hd__decap_12_273 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_295 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_284 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_6_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_ef_sc_hd__decap_12_14 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_25 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_36 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_69 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_58 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_47 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_1_39 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_39/X tt08_integration_0/div_out1_3
+ sky130_fd_sc_hd__mux2_1_39/S sky130_fd_sc_hd__buf_2_7/X sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_17/X sky130_fd_sc_hd__mux2_1_40/A1
+ sky130_fd_sc_hd__nor4b_2_0/Y tt08_integration_0/div_fb3_2 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_28 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_28/X sky130_fd_sc_hd__buf_2_7/X
+ sky130_fd_sc_hd__mux2_1_29/S tt08_integration_0/div_out1_2 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__clkbuf_1_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_16/X uio_in[0]
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__conb_1_16 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_12/A sky130_fd_sc_hd__conb_1_16/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_35 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_24 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__dlymetal6s2s_1_1 VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_1_7/A
+ sky130_fd_sc_hd__clkbuf_1_3/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_fd_sc_hd__nor4b_2_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__buf_2_0/X
+ sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__mux2_1_9/S sky130_fd_sc_hd__buf_2_3/X
+ sky130_fd_sc_hd__nor4b_2
Xsky130_ef_sc_hd__decap_12_296 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_263 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_285 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_274 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_252 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_ef_sc_hd__decap_12_241 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_230 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_6_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_ef_sc_hd__decap_12_26 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_15 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_37 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_59 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_48 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_1_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_18/X sky130_fd_sc_hd__mux2_1_8/A1
+ sky130_fd_sc_hd__mux2_1_23/S tt08_integration_0/div_fb2_3 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__mux2_1_29 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_29/X sky130_fd_sc_hd__mux2_1_4/A1
+ sky130_fd_sc_hd__mux2_1_29/S tt08_integration_0/div_out3_2 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_4_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkbuf_1_17 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_5/A ui_in[4]
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__conb_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_0/A sky130_fd_sc_hd__conb_1_0/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_17 VGND VPWR VGND VPWR uio_oe[0] sky130_fd_sc_hd__conb_1_17/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_36 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_25 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_14 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__dlymetal6s2s_1_2 VPWR VGND VGND VPWR sky130_fd_sc_hd__dfstp_1_2/SET_B
+ sky130_fd_sc_hd__clkbuf_2_1/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_ef_sc_hd__decap_12_297 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_286 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_253 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_275 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_264 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_ef_sc_hd__decap_12_220 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_242 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_231 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_6_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_ef_sc_hd__decap_12_27 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_38 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_16 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_49 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__nor4bb_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__nor4bb_1_0/A sky130_fd_sc_hd__mux2_1_37/S
+ sky130_fd_sc_hd__buf_2_9/A sky130_fd_sc_hd__nand4b_1_0/B sky130_fd_sc_hd__buf_2_8/A
+ sky130_fd_sc_hd__nor4bb_1
Xsky130_fd_sc_hd__mux2_1_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_19/X sky130_fd_sc_hd__buf_2_7/A
+ sky130_fd_sc_hd__mux2_1_23/S tt08_integration_0/div_fb1_3 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_4_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkbuf_1_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_4/A ui_in[7]
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__conb_1_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_2/A sky130_fd_sc_hd__conb_1_1/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__conb_1_18 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_16/A sky130_fd_sc_hd__conb_1_18/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_26 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_37 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_15 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__dlymetal6s2s_1_3 VPWR VGND VGND VPWR sky130_fd_sc_hd__dfstp_1_11/SET_B
+ sky130_fd_sc_hd__clkbuf_2_0/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_ef_sc_hd__decap_12_210 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_276 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_265 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_287 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_298 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_254 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_ef_sc_hd__decap_12_243 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_221 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_232 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_6_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_ef_sc_hd__decap_12_17 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_39 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_28 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__clkbuf_1_19 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_37/A1 sky130_fd_sc_hd__buf_2_7/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__conb_1_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_1/A sky130_fd_sc_hd__conb_1_2/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux4_2_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux4_2_0/S0 sky130_fd_sc_hd__buf_4_19/A
+ sky130_fd_sc_hd__buf_4_17/A sky130_fd_sc_hd__mux4_2_0/S1 sky130_fd_sc_hd__buf_4_20/A
+ sky130_fd_sc_hd__mux4_2_3/A0 sky130_fd_sc_hd__mux4_2_0/X sky130_fd_sc_hd__mux4_2
Xsky130_fd_sc_hd__decap_8_27 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_38 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_16 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__dlymetal6s2s_1_4 VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_2_2/A
+ sky130_fd_sc_hd__clkbuf_1_1/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_ef_sc_hd__decap_12_200 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_244 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_222 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_233 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_211 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_299 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_266 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_277 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_255 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_288 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_8_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_6_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_ef_sc_hd__decap_12_18 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_29 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_4_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__mux4_2_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux4_2_1/S0 sky130_fd_sc_hd__buf_4_20/A
+ sky130_fd_sc_hd__buf_4_17/A sky130_fd_sc_hd__mux4_2_1/S1 sky130_fd_sc_hd__buf_4_18/A
+ sky130_fd_sc_hd__mux4_2_2/A0 sky130_fd_sc_hd__mux4_2_1/X sky130_fd_sc_hd__mux4_2
Xsky130_fd_sc_hd__conb_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_3/A sky130_fd_sc_hd__conb_1_3/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_8_28 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_39 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_17 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__dlymetal6s2s_1_5 VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_1_3/A
+ sky130_fd_sc_hd__clkbuf_1_11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_ef_sc_hd__decap_12_278 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_267 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_256 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_201 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_245 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_212 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_234 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_223 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_289 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_6_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_ef_sc_hd__decap_12_19 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_6_50 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkbuf_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_0/X sky130_fd_sc_hd__clkbuf_1_9/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_4_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_13/A sky130_fd_sc_hd__conb_1_4/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__mux4_2_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux4_2_2/S0 sky130_fd_sc_hd__buf_4_19/A
+ sky130_fd_sc_hd__buf_4_17/A sky130_fd_sc_hd__mux4_2_2/S1 sky130_fd_sc_hd__buf_4_18/A
+ sky130_fd_sc_hd__mux4_2_2/A0 sky130_fd_sc_hd__mux4_2_2/X sky130_fd_sc_hd__mux4_2
Xsky130_fd_sc_hd__decap_8_29 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__decap_8_18 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__dlymetal6s2s_1_6 VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_1_10/A
+ sky130_fd_sc_hd__clkbuf_1_11/X sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_ef_sc_hd__decap_12_268 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_279 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_257 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_202 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_224 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_246 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_213 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_235 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_6_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_51 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_40 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkbuf_1_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_1/A sky130_fd_sc_hd__clkbuf_1_1/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_4_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__mux4_2_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux4_2_3/S0 sky130_fd_sc_hd__buf_4_20/A
+ sky130_fd_sc_hd__buf_4_19/A sky130_fd_sc_hd__mux4_2_3/S1 sky130_fd_sc_hd__buf_4_18/A
+ sky130_fd_sc_hd__mux4_2_3/A0 sky130_fd_sc_hd__mux4_2_3/X sky130_fd_sc_hd__mux4_2
Xsky130_fd_sc_hd__conb_1_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_11/A sky130_fd_sc_hd__conb_1_5/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_3_30 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__clkbuf_2_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_10/A sky130_fd_sc_hd__dfstp_1_9/CLK
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__decap_8_19 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_8
Xsky130_fd_sc_hd__dlymetal6s2s_1_7 VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_1_1/A
+ sky130_fd_sc_hd__dlymetal6s2s_1_7/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_ef_sc_hd__decap_12_269 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_258 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_203 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_236 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_214 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_247 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_225 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_6_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_30 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_41 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_52 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkbuf_1_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_5/A sky130_fd_sc_hd__clkbuf_2_2/X
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_4_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_6/A sky130_fd_sc_hd__conb_1_6/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_3_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_31 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__clkbuf_2_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_5/A sky130_fd_sc_hd__nor4bb_1_0/A
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__dlymetal6s2s_1_8 VPWR VGND VGND VPWR sky130_fd_sc_hd__clkbuf_2_10/A
+ sky130_fd_sc_hd__clkbuf_1_10/A sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_ef_sc_hd__decap_12_204 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_215 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_226 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_259 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_248 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_237 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__decap_6_42 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_31 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_53 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_20 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkbuf_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_5/A sky130_fd_sc_hd__clkbuf_1_3/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_4_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_7 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_14/A sky130_fd_sc_hd__conb_1_7/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_3_21 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__clkbuf_2_12 VGND VPWR VGND VPWR sky130_fd_sc_hd__nor4bb_1_0/A sky130_fd_sc_hd__nor4b_4_0/A
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__dlymetal6s2s_1_9 VPWR VGND VGND VPWR sky130_fd_sc_hd__dfstp_1_10/CLK
+ sky130_fd_sc_hd__dfstp_1_9/CLK sky130_fd_sc_hd__dlymetal6s2s_1
Xsky130_fd_sc_hd__dfrtp_1_30 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_7/A sky130_fd_sc_hd__mux2_1_43/X
+ sky130_fd_sc_hd__clkbuf_2_2/A sky130_fd_sc_hd__mux4_2_2/S0 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_205 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_216 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_249 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_238 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_227 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__nor4_4_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_5/X sky130_fd_sc_hd__buf_2_3/X
+ sky130_fd_sc_hd__nor4_4_0/Y sky130_fd_sc_hd__buf_2_4/X sky130_fd_sc_hd__buf_2_0/X
+ sky130_fd_sc_hd__nor4_4
Xsky130_fd_sc_hd__mux2_1_0 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_0/X sky130_fd_sc_hd__buf_2_7/X
+ sky130_fd_sc_hd__mux2_1_5/S sky130_fd_sc_hd__mux2_1_0/A0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_6_43 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_54 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_32 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_10 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_21 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkbuf_1_4 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_4/X sky130_fd_sc_hd__clkbuf_1_6/X
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_4_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_8 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_15/A sky130_fd_sc_hd__conb_1_8/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_3_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_33 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__clkbuf_2_13 VGND VPWR VGND VPWR ui_in[3] sky130_fd_sc_hd__clkbuf_2_3/A
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__dfrtp_1_20 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_10/A sky130_fd_sc_hd__mux2_1_31/X
+ sky130_fd_sc_hd__clkbuf_2_8/A sky130_fd_sc_hd__mux4_2_1/S1 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfrtp_1_31 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_7/A sky130_fd_sc_hd__mux2_1_42/X
+ sky130_fd_sc_hd__clkbuf_2_2/A sky130_fd_sc_hd__mux4_2_2/S1 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_206 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_239 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_217 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_228 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_1_1 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_1/X sky130_fd_sc_hd__mux2_1_3/A1
+ sky130_fd_sc_hd__mux2_1_5/S sky130_fd_sc_hd__mux2_1_1/A0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_6_44 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_33 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_11 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_22 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_55 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkbuf_1_5 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_5/X sky130_fd_sc_hd__clkbuf_1_5/A
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_4_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__decap_4
Xsky130_fd_sc_hd__conb_1_9 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_4_10/A sky130_fd_sc_hd__conb_1_9/HI
+ sky130_fd_sc_hd__conb_1
Xsky130_fd_sc_hd__decap_3_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__clkbuf_2_14 VGND VPWR VGND VPWR ui_in[2] sky130_fd_sc_hd__clkbuf_2_9/A
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__dfrtp_1_21 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_10/A sky130_fd_sc_hd__mux2_1_30/X
+ sky130_fd_sc_hd__clkbuf_2_8/A sky130_fd_sc_hd__mux4_2_1/S0 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfrtp_1_10 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__mux2_1_20/X
+ sky130_fd_sc_hd__clkbuf_2_2/X tt08_integration_0/div_fb3_3 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_229 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_207 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_218 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xtt08_integration_0 tt08_integration_0/div_fb0_1 tt08_integration_0/div_fb1_1 tt08_integration_0/div_fb2_1
+ tt08_integration_0/div_fb3_1 tt08_integration_0/div_out0_1 sky130_fd_sc_hd__mux2_1_3/A0
+ sky130_fd_sc_hd__dfrtp_1_4/Q tt08_integration_0/div_out3_1 tt08_integration_0/div_out3_2
+ tt08_integration_0/div_out1_2 tt08_integration_0/div_out2_2 sky130_fd_sc_hd__dfstp_1_9/Q
+ tt08_integration_0/div_fb3_2 tt08_integration_0/div_fb2_2 tt08_integration_0/div_fb1_2
+ tt08_integration_0/div_fb0_2 tt08_integration_0/div_out3_3 tt08_integration_0/div_out1_3
+ tt08_integration_0/div_out2_3 tt08_integration_0/div_out0_3 tt08_integration_0/div_fb3_3
+ tt08_integration_0/div_fb2_3 tt08_integration_0/div_fb1_3 tt08_integration_0/div_fb0_3
+ tt08_integration_0/div_fb0_0 tt08_integration_0/div_fb1_0 tt08_integration_0/div_fb2_0
+ tt08_integration_0/div_fb3_0 sky130_fd_sc_hd__mux2_1_5/A0 sky130_fd_sc_hd__mux2_1_1/A0
+ sky130_fd_sc_hd__mux2_1_0/A0 sky130_fd_sc_hd__mux2_1_4/A0 tt08_integration_0/enb_0
+ sky130_fd_sc_hd__mux4_2_0/X VPWR VPWR sky130_fd_sc_hd__dfstp_1_2/Q VGND VPWR VGND
+ VPWR sky130_fd_sc_hd__mux4_2_2/X sky130_fd_sc_hd__clkbuf_1_12/A VGND sky130_fd_sc_hd__buf_4_20/A
+ VGND VPWR sky130_fd_sc_hd__buf_4_19/A VPWR VGND VPWR sky130_fd_sc_hd__buf_4_18/A
+ VPWR VPWR VPWR VPWR VGND VPWR sky130_fd_sc_hd__mux4_2_1/X VPWR VGND sky130_fd_sc_hd__mux4_2_3/X
+ VGND VPWR sky130_fd_sc_hd__dfstp_1_6/Q sky130_fd_sc_hd__buf_4_17/A sky130_fd_sc_hd__dfstp_1_8/Q
+ VPWR VGND VGND VGND VGND VGND tt08_integration
Xsky130_fd_sc_hd__mux2_1_2 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_2/X sky130_fd_sc_hd__buf_2_6/X
+ sky130_fd_sc_hd__mux2_1_2/S tt08_integration_0/enb_0 sky130_fd_sc_hd__mux2_1
Xsky130_fd_sc_hd__decap_6_12 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_23 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_34 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_45 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__decap_6_56 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_6
Xsky130_fd_sc_hd__clkbuf_1_6 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_6/X sky130_fd_sc_hd__clkbuf_1_7/X
+ sky130_fd_sc_hd__clkbuf_1
Xsky130_fd_sc_hd__decap_3_24 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_35 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__decap_3_13 VPWR VGND VGND VPWR sky130_fd_sc_hd__decap_3
Xsky130_fd_sc_hd__clkbuf_2_15 VGND VPWR VGND VPWR sky130_fd_sc_hd__buf_2_6/A sky130_fd_sc_hd__mux2_1_35/A1
+ sky130_fd_sc_hd__clkbuf_2
Xsky130_fd_sc_hd__dfrtp_1_22 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_2_10/A sky130_fd_sc_hd__mux2_1_32/X
+ sky130_fd_sc_hd__clkbuf_2_8/A sky130_fd_sc_hd__mux4_2_0/S1 sky130_fd_sc_hd__dfrtp_1
Xsky130_fd_sc_hd__dfrtp_1_11 VGND VPWR VGND VPWR sky130_fd_sc_hd__clkbuf_1_7/X sky130_fd_sc_hd__mux2_1_18/X
+ sky130_fd_sc_hd__clkbuf_2_2/X tt08_integration_0/div_fb2_3 sky130_fd_sc_hd__dfrtp_1
Xsky130_ef_sc_hd__decap_12_208 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_ef_sc_hd__decap_12_219 VGND VPWR VGND VPWR sky130_ef_sc_hd__decap_12
Xsky130_fd_sc_hd__mux2_1_3 VGND VPWR VGND VPWR sky130_fd_sc_hd__mux2_1_3/X sky130_fd_sc_hd__mux2_1_3/A1
+ sky130_fd_sc_hd__mux2_1_3/S sky130_fd_sc_hd__mux2_1_3/A0 sky130_fd_sc_hd__mux2_1
.ends

